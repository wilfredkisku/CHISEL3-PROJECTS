module BufferMemorySystem(
  input        clock,
  input        reset,
  input        io_enable,
  input        io_write,
  input  [3:0] io_addr,
  input  [7:0] io_adcValues_0,
  input  [7:0] io_adcValues_1,
  input  [7:0] io_adcValues_2,
  input  [7:0] io_adcValues_3,
  input  [7:0] io_adcValues_4,
  input  [7:0] io_adcValues_5,
  input  [7:0] io_adcValues_6,
  input  [7:0] io_adcValues_7,
  input  [7:0] io_adcValues_8,
  input  [7:0] io_adcValues_9,
  input  [7:0] io_adcValues_10,
  input  [7:0] io_adcValues_11,
  input  [7:0] io_adcValues_12,
  input  [7:0] io_adcValues_13,
  input  [7:0] io_adcValues_14,
  input  [7:0] io_adcValues_15,
  input  [7:0] io_adcValues_16,
  input  [7:0] io_adcValues_17,
  input  [7:0] io_adcValues_18,
  input  [7:0] io_adcValues_19,
  input  [7:0] io_adcValues_20,
  input  [7:0] io_adcValues_21,
  input  [7:0] io_adcValues_22,
  input  [7:0] io_adcValues_23,
  input  [7:0] io_adcValues_24,
  input  [7:0] io_adcValues_25,
  input  [7:0] io_adcValues_26,
  input  [7:0] io_adcValues_27,
  input  [7:0] io_adcValues_28,
  input  [7:0] io_adcValues_29,
  input  [7:0] io_adcValues_30,
  input  [7:0] io_adcValues_31,
  input  [7:0] io_adcValues_32,
  input  [7:0] io_adcValues_33,
  input  [7:0] io_adcValues_34,
  input  [7:0] io_adcValues_35,
  input  [7:0] io_adcValues_36,
  input  [7:0] io_adcValues_37,
  input  [7:0] io_adcValues_38,
  input  [7:0] io_adcValues_39,
  input  [7:0] io_adcValues_40,
  input  [7:0] io_adcValues_41,
  input  [7:0] io_adcValues_42,
  input  [7:0] io_adcValues_43,
  input  [7:0] io_adcValues_44,
  input  [7:0] io_adcValues_45,
  input  [7:0] io_adcValues_46,
  input  [7:0] io_adcValues_47,
  input  [7:0] io_adcValues_48,
  input  [7:0] io_adcValues_49,
  input  [7:0] io_adcValues_50,
  input  [7:0] io_adcValues_51,
  input  [7:0] io_adcValues_52,
  input  [7:0] io_adcValues_53,
  input  [7:0] io_adcValues_54,
  input  [7:0] io_adcValues_55,
  input  [7:0] io_adcValues_56,
  input  [7:0] io_adcValues_57,
  input  [7:0] io_adcValues_58,
  input  [7:0] io_adcValues_59,
  input  [7:0] io_adcValues_60,
  input  [7:0] io_adcValues_61,
  input  [7:0] io_adcValues_62,
  input  [7:0] io_adcValues_63,
  input  [7:0] io_adcValues_64,
  input  [7:0] io_adcValues_65,
  input  [7:0] io_adcValues_66,
  input  [7:0] io_adcValues_67,
  input  [7:0] io_adcValues_68,
  input  [7:0] io_adcValues_69,
  input  [7:0] io_adcValues_70,
  input  [7:0] io_adcValues_71,
  input  [7:0] io_adcValues_72,
  input  [7:0] io_adcValues_73,
  input  [7:0] io_adcValues_74,
  input  [7:0] io_adcValues_75,
  input  [7:0] io_adcValues_76,
  input  [7:0] io_adcValues_77,
  input  [7:0] io_adcValues_78,
  input  [7:0] io_adcValues_79,
  input  [7:0] io_adcValues_80,
  input  [7:0] io_adcValues_81,
  input  [7:0] io_adcValues_82,
  input  [7:0] io_adcValues_83,
  input  [7:0] io_adcValues_84,
  input  [7:0] io_adcValues_85,
  input  [7:0] io_adcValues_86,
  input  [7:0] io_adcValues_87,
  input  [7:0] io_adcValues_88,
  input  [7:0] io_adcValues_89,
  input  [7:0] io_adcValues_90,
  input  [7:0] io_adcValues_91,
  input  [7:0] io_adcValues_92,
  input  [7:0] io_adcValues_93,
  input  [7:0] io_adcValues_94,
  input  [7:0] io_adcValues_95,
  input  [7:0] io_adcValues_96,
  input  [7:0] io_adcValues_97,
  input  [7:0] io_adcValues_98,
  input  [7:0] io_adcValues_99,
  input  [7:0] io_adcValues_100,
  input  [7:0] io_adcValues_101,
  input  [7:0] io_adcValues_102,
  input  [7:0] io_adcValues_103,
  input  [7:0] io_adcValues_104,
  input  [7:0] io_adcValues_105,
  input  [7:0] io_adcValues_106,
  input  [7:0] io_adcValues_107,
  input  [7:0] io_adcValues_108,
  input  [7:0] io_adcValues_109,
  input  [7:0] io_adcValues_110,
  input  [7:0] io_adcValues_111,
  input  [7:0] io_adcValues_112,
  input  [7:0] io_adcValues_113,
  input  [7:0] io_adcValues_114,
  input  [7:0] io_adcValues_115,
  input  [7:0] io_adcValues_116,
  input  [7:0] io_adcValues_117,
  input  [7:0] io_adcValues_118,
  input  [7:0] io_adcValues_119,
  input  [7:0] io_adcValues_120,
  input  [7:0] io_adcValues_121,
  input  [7:0] io_adcValues_122,
  input  [7:0] io_adcValues_123,
  input  [7:0] io_adcValues_124,
  input  [7:0] io_adcValues_125,
  input  [7:0] io_adcValues_126,
  input  [7:0] io_adcValues_127,
  output [7:0] io_dataOut_0,
  output [7:0] io_dataOut_1,
  output [7:0] io_dataOut_2,
  output [7:0] io_dataOut_3,
  output [7:0] io_dataOut_4,
  output [7:0] io_dataOut_5,
  output [7:0] io_dataOut_6,
  output [7:0] io_dataOut_7,
  output [7:0] io_dataOut_8,
  output [7:0] io_dataOut_9,
  output [7:0] io_dataOut_10,
  output [7:0] io_dataOut_11,
  output [7:0] io_dataOut_12,
  output [7:0] io_dataOut_13,
  output [7:0] io_dataOut_14,
  output [7:0] io_dataOut_15,
  output [7:0] io_dataOut_16,
  output [7:0] io_dataOut_17,
  output [7:0] io_dataOut_18,
  output [7:0] io_dataOut_19,
  output [7:0] io_dataOut_20,
  output [7:0] io_dataOut_21,
  output [7:0] io_dataOut_22,
  output [7:0] io_dataOut_23,
  output [7:0] io_dataOut_24,
  output [7:0] io_dataOut_25,
  output [7:0] io_dataOut_26,
  output [7:0] io_dataOut_27,
  output [7:0] io_dataOut_28,
  output [7:0] io_dataOut_29,
  output [7:0] io_dataOut_30,
  output [7:0] io_dataOut_31,
  output [7:0] io_dataOut_32,
  output [7:0] io_dataOut_33,
  output [7:0] io_dataOut_34,
  output [7:0] io_dataOut_35,
  output [7:0] io_dataOut_36,
  output [7:0] io_dataOut_37,
  output [7:0] io_dataOut_38,
  output [7:0] io_dataOut_39,
  output [7:0] io_dataOut_40,
  output [7:0] io_dataOut_41,
  output [7:0] io_dataOut_42,
  output [7:0] io_dataOut_43,
  output [7:0] io_dataOut_44,
  output [7:0] io_dataOut_45,
  output [7:0] io_dataOut_46,
  output [7:0] io_dataOut_47,
  output [7:0] io_dataOut_48,
  output [7:0] io_dataOut_49,
  output [7:0] io_dataOut_50,
  output [7:0] io_dataOut_51,
  output [7:0] io_dataOut_52,
  output [7:0] io_dataOut_53,
  output [7:0] io_dataOut_54,
  output [7:0] io_dataOut_55,
  output [7:0] io_dataOut_56,
  output [7:0] io_dataOut_57,
  output [7:0] io_dataOut_58,
  output [7:0] io_dataOut_59,
  output [7:0] io_dataOut_60,
  output [7:0] io_dataOut_61,
  output [7:0] io_dataOut_62,
  output [7:0] io_dataOut_63,
  output [7:0] io_dataOut_64,
  output [7:0] io_dataOut_65,
  output [7:0] io_dataOut_66,
  output [7:0] io_dataOut_67,
  output [7:0] io_dataOut_68,
  output [7:0] io_dataOut_69,
  output [7:0] io_dataOut_70,
  output [7:0] io_dataOut_71,
  output [7:0] io_dataOut_72,
  output [7:0] io_dataOut_73,
  output [7:0] io_dataOut_74,
  output [7:0] io_dataOut_75,
  output [7:0] io_dataOut_76,
  output [7:0] io_dataOut_77,
  output [7:0] io_dataOut_78,
  output [7:0] io_dataOut_79,
  output [7:0] io_dataOut_80,
  output [7:0] io_dataOut_81,
  output [7:0] io_dataOut_82,
  output [7:0] io_dataOut_83,
  output [7:0] io_dataOut_84,
  output [7:0] io_dataOut_85,
  output [7:0] io_dataOut_86,
  output [7:0] io_dataOut_87,
  output [7:0] io_dataOut_88,
  output [7:0] io_dataOut_89,
  output [7:0] io_dataOut_90,
  output [7:0] io_dataOut_91,
  output [7:0] io_dataOut_92,
  output [7:0] io_dataOut_93,
  output [7:0] io_dataOut_94,
  output [7:0] io_dataOut_95,
  output [7:0] io_dataOut_96,
  output [7:0] io_dataOut_97,
  output [7:0] io_dataOut_98,
  output [7:0] io_dataOut_99,
  output [7:0] io_dataOut_100,
  output [7:0] io_dataOut_101,
  output [7:0] io_dataOut_102,
  output [7:0] io_dataOut_103,
  output [7:0] io_dataOut_104,
  output [7:0] io_dataOut_105,
  output [7:0] io_dataOut_106,
  output [7:0] io_dataOut_107,
  output [7:0] io_dataOut_108,
  output [7:0] io_dataOut_109,
  output [7:0] io_dataOut_110,
  output [7:0] io_dataOut_111,
  output [7:0] io_dataOut_112,
  output [7:0] io_dataOut_113,
  output [7:0] io_dataOut_114,
  output [7:0] io_dataOut_115,
  output [7:0] io_dataOut_116,
  output [7:0] io_dataOut_117,
  output [7:0] io_dataOut_118,
  output [7:0] io_dataOut_119,
  output [7:0] io_dataOut_120,
  output [7:0] io_dataOut_121,
  output [7:0] io_dataOut_122,
  output [7:0] io_dataOut_123,
  output [7:0] io_dataOut_124,
  output [7:0] io_dataOut_125,
  output [7:0] io_dataOut_126,
  output [7:0] io_dataOut_127
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_381;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] mem_0 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_0_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_0_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_0_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_0_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_0_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_0_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_0_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_0_MPORT_1_en_pipe_0;
  reg [3:0] mem_0_MPORT_1_addr_pipe_0;
  reg [7:0] mem_1 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_1_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_1_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_1_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_1_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_1_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_1_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_1_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_1_MPORT_1_en_pipe_0;
  reg [3:0] mem_1_MPORT_1_addr_pipe_0;
  reg [7:0] mem_2 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_2_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_2_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_2_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_2_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_2_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_2_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_2_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_2_MPORT_1_en_pipe_0;
  reg [3:0] mem_2_MPORT_1_addr_pipe_0;
  reg [7:0] mem_3 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_3_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_3_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_3_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_3_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_3_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_3_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_3_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_3_MPORT_1_en_pipe_0;
  reg [3:0] mem_3_MPORT_1_addr_pipe_0;
  reg [7:0] mem_4 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_4_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_4_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_4_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_4_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_4_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_4_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_4_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_4_MPORT_1_en_pipe_0;
  reg [3:0] mem_4_MPORT_1_addr_pipe_0;
  reg [7:0] mem_5 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_5_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_5_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_5_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_5_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_5_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_5_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_5_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_5_MPORT_1_en_pipe_0;
  reg [3:0] mem_5_MPORT_1_addr_pipe_0;
  reg [7:0] mem_6 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_6_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_6_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_6_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_6_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_6_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_6_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_6_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_6_MPORT_1_en_pipe_0;
  reg [3:0] mem_6_MPORT_1_addr_pipe_0;
  reg [7:0] mem_7 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_7_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_7_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_7_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_7_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_7_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_7_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_7_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_7_MPORT_1_en_pipe_0;
  reg [3:0] mem_7_MPORT_1_addr_pipe_0;
  reg [7:0] mem_8 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_8_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_8_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_8_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_8_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_8_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_8_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_8_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_8_MPORT_1_en_pipe_0;
  reg [3:0] mem_8_MPORT_1_addr_pipe_0;
  reg [7:0] mem_9 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_9_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_9_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_9_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_9_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_9_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_9_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_9_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_9_MPORT_1_en_pipe_0;
  reg [3:0] mem_9_MPORT_1_addr_pipe_0;
  reg [7:0] mem_10 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_10_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_10_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_10_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_10_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_10_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_10_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_10_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_10_MPORT_1_en_pipe_0;
  reg [3:0] mem_10_MPORT_1_addr_pipe_0;
  reg [7:0] mem_11 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_11_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_11_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_11_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_11_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_11_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_11_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_11_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_11_MPORT_1_en_pipe_0;
  reg [3:0] mem_11_MPORT_1_addr_pipe_0;
  reg [7:0] mem_12 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_12_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_12_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_12_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_12_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_12_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_12_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_12_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_12_MPORT_1_en_pipe_0;
  reg [3:0] mem_12_MPORT_1_addr_pipe_0;
  reg [7:0] mem_13 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_13_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_13_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_13_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_13_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_13_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_13_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_13_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_13_MPORT_1_en_pipe_0;
  reg [3:0] mem_13_MPORT_1_addr_pipe_0;
  reg [7:0] mem_14 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_14_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_14_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_14_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_14_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_14_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_14_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_14_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_14_MPORT_1_en_pipe_0;
  reg [3:0] mem_14_MPORT_1_addr_pipe_0;
  reg [7:0] mem_15 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_15_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_15_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_15_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_15_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_15_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_15_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_15_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_15_MPORT_1_en_pipe_0;
  reg [3:0] mem_15_MPORT_1_addr_pipe_0;
  reg [7:0] mem_16 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_16_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_16_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_16_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_16_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_16_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_16_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_16_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_16_MPORT_1_en_pipe_0;
  reg [3:0] mem_16_MPORT_1_addr_pipe_0;
  reg [7:0] mem_17 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_17_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_17_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_17_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_17_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_17_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_17_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_17_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_17_MPORT_1_en_pipe_0;
  reg [3:0] mem_17_MPORT_1_addr_pipe_0;
  reg [7:0] mem_18 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_18_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_18_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_18_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_18_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_18_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_18_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_18_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_18_MPORT_1_en_pipe_0;
  reg [3:0] mem_18_MPORT_1_addr_pipe_0;
  reg [7:0] mem_19 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_19_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_19_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_19_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_19_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_19_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_19_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_19_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_19_MPORT_1_en_pipe_0;
  reg [3:0] mem_19_MPORT_1_addr_pipe_0;
  reg [7:0] mem_20 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_20_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_20_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_20_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_20_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_20_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_20_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_20_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_20_MPORT_1_en_pipe_0;
  reg [3:0] mem_20_MPORT_1_addr_pipe_0;
  reg [7:0] mem_21 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_21_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_21_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_21_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_21_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_21_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_21_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_21_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_21_MPORT_1_en_pipe_0;
  reg [3:0] mem_21_MPORT_1_addr_pipe_0;
  reg [7:0] mem_22 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_22_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_22_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_22_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_22_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_22_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_22_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_22_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_22_MPORT_1_en_pipe_0;
  reg [3:0] mem_22_MPORT_1_addr_pipe_0;
  reg [7:0] mem_23 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_23_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_23_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_23_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_23_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_23_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_23_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_23_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_23_MPORT_1_en_pipe_0;
  reg [3:0] mem_23_MPORT_1_addr_pipe_0;
  reg [7:0] mem_24 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_24_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_24_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_24_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_24_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_24_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_24_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_24_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_24_MPORT_1_en_pipe_0;
  reg [3:0] mem_24_MPORT_1_addr_pipe_0;
  reg [7:0] mem_25 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_25_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_25_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_25_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_25_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_25_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_25_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_25_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_25_MPORT_1_en_pipe_0;
  reg [3:0] mem_25_MPORT_1_addr_pipe_0;
  reg [7:0] mem_26 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_26_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_26_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_26_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_26_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_26_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_26_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_26_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_26_MPORT_1_en_pipe_0;
  reg [3:0] mem_26_MPORT_1_addr_pipe_0;
  reg [7:0] mem_27 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_27_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_27_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_27_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_27_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_27_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_27_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_27_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_27_MPORT_1_en_pipe_0;
  reg [3:0] mem_27_MPORT_1_addr_pipe_0;
  reg [7:0] mem_28 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_28_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_28_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_28_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_28_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_28_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_28_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_28_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_28_MPORT_1_en_pipe_0;
  reg [3:0] mem_28_MPORT_1_addr_pipe_0;
  reg [7:0] mem_29 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_29_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_29_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_29_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_29_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_29_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_29_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_29_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_29_MPORT_1_en_pipe_0;
  reg [3:0] mem_29_MPORT_1_addr_pipe_0;
  reg [7:0] mem_30 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_30_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_30_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_30_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_30_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_30_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_30_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_30_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_30_MPORT_1_en_pipe_0;
  reg [3:0] mem_30_MPORT_1_addr_pipe_0;
  reg [7:0] mem_31 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_31_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_31_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_31_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_31_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_31_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_31_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_31_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_31_MPORT_1_en_pipe_0;
  reg [3:0] mem_31_MPORT_1_addr_pipe_0;
  reg [7:0] mem_32 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_32_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_32_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_32_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_32_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_32_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_32_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_32_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_32_MPORT_1_en_pipe_0;
  reg [3:0] mem_32_MPORT_1_addr_pipe_0;
  reg [7:0] mem_33 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_33_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_33_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_33_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_33_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_33_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_33_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_33_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_33_MPORT_1_en_pipe_0;
  reg [3:0] mem_33_MPORT_1_addr_pipe_0;
  reg [7:0] mem_34 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_34_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_34_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_34_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_34_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_34_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_34_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_34_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_34_MPORT_1_en_pipe_0;
  reg [3:0] mem_34_MPORT_1_addr_pipe_0;
  reg [7:0] mem_35 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_35_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_35_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_35_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_35_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_35_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_35_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_35_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_35_MPORT_1_en_pipe_0;
  reg [3:0] mem_35_MPORT_1_addr_pipe_0;
  reg [7:0] mem_36 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_36_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_36_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_36_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_36_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_36_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_36_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_36_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_36_MPORT_1_en_pipe_0;
  reg [3:0] mem_36_MPORT_1_addr_pipe_0;
  reg [7:0] mem_37 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_37_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_37_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_37_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_37_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_37_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_37_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_37_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_37_MPORT_1_en_pipe_0;
  reg [3:0] mem_37_MPORT_1_addr_pipe_0;
  reg [7:0] mem_38 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_38_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_38_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_38_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_38_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_38_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_38_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_38_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_38_MPORT_1_en_pipe_0;
  reg [3:0] mem_38_MPORT_1_addr_pipe_0;
  reg [7:0] mem_39 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_39_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_39_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_39_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_39_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_39_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_39_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_39_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_39_MPORT_1_en_pipe_0;
  reg [3:0] mem_39_MPORT_1_addr_pipe_0;
  reg [7:0] mem_40 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_40_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_40_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_40_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_40_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_40_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_40_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_40_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_40_MPORT_1_en_pipe_0;
  reg [3:0] mem_40_MPORT_1_addr_pipe_0;
  reg [7:0] mem_41 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_41_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_41_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_41_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_41_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_41_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_41_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_41_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_41_MPORT_1_en_pipe_0;
  reg [3:0] mem_41_MPORT_1_addr_pipe_0;
  reg [7:0] mem_42 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_42_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_42_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_42_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_42_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_42_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_42_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_42_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_42_MPORT_1_en_pipe_0;
  reg [3:0] mem_42_MPORT_1_addr_pipe_0;
  reg [7:0] mem_43 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_43_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_43_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_43_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_43_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_43_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_43_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_43_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_43_MPORT_1_en_pipe_0;
  reg [3:0] mem_43_MPORT_1_addr_pipe_0;
  reg [7:0] mem_44 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_44_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_44_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_44_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_44_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_44_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_44_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_44_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_44_MPORT_1_en_pipe_0;
  reg [3:0] mem_44_MPORT_1_addr_pipe_0;
  reg [7:0] mem_45 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_45_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_45_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_45_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_45_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_45_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_45_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_45_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_45_MPORT_1_en_pipe_0;
  reg [3:0] mem_45_MPORT_1_addr_pipe_0;
  reg [7:0] mem_46 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_46_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_46_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_46_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_46_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_46_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_46_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_46_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_46_MPORT_1_en_pipe_0;
  reg [3:0] mem_46_MPORT_1_addr_pipe_0;
  reg [7:0] mem_47 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_47_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_47_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_47_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_47_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_47_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_47_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_47_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_47_MPORT_1_en_pipe_0;
  reg [3:0] mem_47_MPORT_1_addr_pipe_0;
  reg [7:0] mem_48 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_48_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_48_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_48_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_48_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_48_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_48_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_48_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_48_MPORT_1_en_pipe_0;
  reg [3:0] mem_48_MPORT_1_addr_pipe_0;
  reg [7:0] mem_49 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_49_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_49_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_49_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_49_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_49_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_49_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_49_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_49_MPORT_1_en_pipe_0;
  reg [3:0] mem_49_MPORT_1_addr_pipe_0;
  reg [7:0] mem_50 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_50_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_50_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_50_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_50_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_50_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_50_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_50_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_50_MPORT_1_en_pipe_0;
  reg [3:0] mem_50_MPORT_1_addr_pipe_0;
  reg [7:0] mem_51 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_51_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_51_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_51_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_51_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_51_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_51_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_51_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_51_MPORT_1_en_pipe_0;
  reg [3:0] mem_51_MPORT_1_addr_pipe_0;
  reg [7:0] mem_52 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_52_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_52_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_52_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_52_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_52_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_52_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_52_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_52_MPORT_1_en_pipe_0;
  reg [3:0] mem_52_MPORT_1_addr_pipe_0;
  reg [7:0] mem_53 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_53_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_53_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_53_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_53_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_53_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_53_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_53_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_53_MPORT_1_en_pipe_0;
  reg [3:0] mem_53_MPORT_1_addr_pipe_0;
  reg [7:0] mem_54 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_54_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_54_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_54_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_54_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_54_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_54_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_54_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_54_MPORT_1_en_pipe_0;
  reg [3:0] mem_54_MPORT_1_addr_pipe_0;
  reg [7:0] mem_55 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_55_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_55_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_55_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_55_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_55_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_55_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_55_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_55_MPORT_1_en_pipe_0;
  reg [3:0] mem_55_MPORT_1_addr_pipe_0;
  reg [7:0] mem_56 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_56_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_56_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_56_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_56_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_56_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_56_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_56_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_56_MPORT_1_en_pipe_0;
  reg [3:0] mem_56_MPORT_1_addr_pipe_0;
  reg [7:0] mem_57 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_57_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_57_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_57_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_57_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_57_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_57_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_57_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_57_MPORT_1_en_pipe_0;
  reg [3:0] mem_57_MPORT_1_addr_pipe_0;
  reg [7:0] mem_58 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_58_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_58_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_58_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_58_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_58_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_58_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_58_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_58_MPORT_1_en_pipe_0;
  reg [3:0] mem_58_MPORT_1_addr_pipe_0;
  reg [7:0] mem_59 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_59_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_59_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_59_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_59_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_59_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_59_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_59_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_59_MPORT_1_en_pipe_0;
  reg [3:0] mem_59_MPORT_1_addr_pipe_0;
  reg [7:0] mem_60 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_60_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_60_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_60_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_60_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_60_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_60_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_60_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_60_MPORT_1_en_pipe_0;
  reg [3:0] mem_60_MPORT_1_addr_pipe_0;
  reg [7:0] mem_61 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_61_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_61_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_61_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_61_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_61_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_61_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_61_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_61_MPORT_1_en_pipe_0;
  reg [3:0] mem_61_MPORT_1_addr_pipe_0;
  reg [7:0] mem_62 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_62_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_62_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_62_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_62_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_62_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_62_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_62_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_62_MPORT_1_en_pipe_0;
  reg [3:0] mem_62_MPORT_1_addr_pipe_0;
  reg [7:0] mem_63 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_63_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_63_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_63_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_63_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_63_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_63_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_63_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_63_MPORT_1_en_pipe_0;
  reg [3:0] mem_63_MPORT_1_addr_pipe_0;
  reg [7:0] mem_64 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_64_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_64_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_64_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_64_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_64_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_64_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_64_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_64_MPORT_1_en_pipe_0;
  reg [3:0] mem_64_MPORT_1_addr_pipe_0;
  reg [7:0] mem_65 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_65_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_65_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_65_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_65_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_65_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_65_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_65_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_65_MPORT_1_en_pipe_0;
  reg [3:0] mem_65_MPORT_1_addr_pipe_0;
  reg [7:0] mem_66 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_66_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_66_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_66_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_66_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_66_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_66_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_66_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_66_MPORT_1_en_pipe_0;
  reg [3:0] mem_66_MPORT_1_addr_pipe_0;
  reg [7:0] mem_67 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_67_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_67_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_67_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_67_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_67_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_67_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_67_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_67_MPORT_1_en_pipe_0;
  reg [3:0] mem_67_MPORT_1_addr_pipe_0;
  reg [7:0] mem_68 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_68_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_68_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_68_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_68_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_68_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_68_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_68_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_68_MPORT_1_en_pipe_0;
  reg [3:0] mem_68_MPORT_1_addr_pipe_0;
  reg [7:0] mem_69 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_69_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_69_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_69_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_69_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_69_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_69_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_69_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_69_MPORT_1_en_pipe_0;
  reg [3:0] mem_69_MPORT_1_addr_pipe_0;
  reg [7:0] mem_70 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_70_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_70_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_70_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_70_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_70_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_70_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_70_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_70_MPORT_1_en_pipe_0;
  reg [3:0] mem_70_MPORT_1_addr_pipe_0;
  reg [7:0] mem_71 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_71_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_71_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_71_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_71_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_71_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_71_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_71_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_71_MPORT_1_en_pipe_0;
  reg [3:0] mem_71_MPORT_1_addr_pipe_0;
  reg [7:0] mem_72 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_72_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_72_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_72_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_72_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_72_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_72_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_72_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_72_MPORT_1_en_pipe_0;
  reg [3:0] mem_72_MPORT_1_addr_pipe_0;
  reg [7:0] mem_73 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_73_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_73_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_73_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_73_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_73_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_73_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_73_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_73_MPORT_1_en_pipe_0;
  reg [3:0] mem_73_MPORT_1_addr_pipe_0;
  reg [7:0] mem_74 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_74_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_74_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_74_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_74_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_74_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_74_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_74_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_74_MPORT_1_en_pipe_0;
  reg [3:0] mem_74_MPORT_1_addr_pipe_0;
  reg [7:0] mem_75 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_75_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_75_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_75_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_75_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_75_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_75_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_75_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_75_MPORT_1_en_pipe_0;
  reg [3:0] mem_75_MPORT_1_addr_pipe_0;
  reg [7:0] mem_76 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_76_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_76_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_76_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_76_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_76_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_76_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_76_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_76_MPORT_1_en_pipe_0;
  reg [3:0] mem_76_MPORT_1_addr_pipe_0;
  reg [7:0] mem_77 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_77_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_77_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_77_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_77_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_77_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_77_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_77_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_77_MPORT_1_en_pipe_0;
  reg [3:0] mem_77_MPORT_1_addr_pipe_0;
  reg [7:0] mem_78 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_78_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_78_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_78_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_78_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_78_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_78_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_78_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_78_MPORT_1_en_pipe_0;
  reg [3:0] mem_78_MPORT_1_addr_pipe_0;
  reg [7:0] mem_79 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_79_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_79_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_79_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_79_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_79_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_79_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_79_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_79_MPORT_1_en_pipe_0;
  reg [3:0] mem_79_MPORT_1_addr_pipe_0;
  reg [7:0] mem_80 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_80_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_80_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_80_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_80_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_80_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_80_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_80_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_80_MPORT_1_en_pipe_0;
  reg [3:0] mem_80_MPORT_1_addr_pipe_0;
  reg [7:0] mem_81 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_81_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_81_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_81_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_81_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_81_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_81_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_81_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_81_MPORT_1_en_pipe_0;
  reg [3:0] mem_81_MPORT_1_addr_pipe_0;
  reg [7:0] mem_82 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_82_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_82_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_82_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_82_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_82_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_82_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_82_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_82_MPORT_1_en_pipe_0;
  reg [3:0] mem_82_MPORT_1_addr_pipe_0;
  reg [7:0] mem_83 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_83_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_83_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_83_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_83_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_83_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_83_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_83_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_83_MPORT_1_en_pipe_0;
  reg [3:0] mem_83_MPORT_1_addr_pipe_0;
  reg [7:0] mem_84 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_84_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_84_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_84_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_84_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_84_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_84_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_84_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_84_MPORT_1_en_pipe_0;
  reg [3:0] mem_84_MPORT_1_addr_pipe_0;
  reg [7:0] mem_85 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_85_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_85_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_85_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_85_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_85_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_85_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_85_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_85_MPORT_1_en_pipe_0;
  reg [3:0] mem_85_MPORT_1_addr_pipe_0;
  reg [7:0] mem_86 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_86_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_86_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_86_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_86_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_86_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_86_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_86_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_86_MPORT_1_en_pipe_0;
  reg [3:0] mem_86_MPORT_1_addr_pipe_0;
  reg [7:0] mem_87 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_87_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_87_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_87_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_87_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_87_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_87_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_87_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_87_MPORT_1_en_pipe_0;
  reg [3:0] mem_87_MPORT_1_addr_pipe_0;
  reg [7:0] mem_88 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_88_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_88_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_88_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_88_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_88_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_88_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_88_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_88_MPORT_1_en_pipe_0;
  reg [3:0] mem_88_MPORT_1_addr_pipe_0;
  reg [7:0] mem_89 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_89_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_89_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_89_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_89_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_89_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_89_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_89_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_89_MPORT_1_en_pipe_0;
  reg [3:0] mem_89_MPORT_1_addr_pipe_0;
  reg [7:0] mem_90 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_90_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_90_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_90_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_90_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_90_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_90_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_90_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_90_MPORT_1_en_pipe_0;
  reg [3:0] mem_90_MPORT_1_addr_pipe_0;
  reg [7:0] mem_91 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_91_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_91_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_91_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_91_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_91_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_91_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_91_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_91_MPORT_1_en_pipe_0;
  reg [3:0] mem_91_MPORT_1_addr_pipe_0;
  reg [7:0] mem_92 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_92_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_92_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_92_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_92_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_92_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_92_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_92_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_92_MPORT_1_en_pipe_0;
  reg [3:0] mem_92_MPORT_1_addr_pipe_0;
  reg [7:0] mem_93 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_93_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_93_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_93_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_93_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_93_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_93_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_93_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_93_MPORT_1_en_pipe_0;
  reg [3:0] mem_93_MPORT_1_addr_pipe_0;
  reg [7:0] mem_94 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_94_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_94_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_94_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_94_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_94_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_94_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_94_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_94_MPORT_1_en_pipe_0;
  reg [3:0] mem_94_MPORT_1_addr_pipe_0;
  reg [7:0] mem_95 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_95_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_95_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_95_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_95_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_95_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_95_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_95_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_95_MPORT_1_en_pipe_0;
  reg [3:0] mem_95_MPORT_1_addr_pipe_0;
  reg [7:0] mem_96 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_96_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_96_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_96_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_96_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_96_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_96_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_96_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_96_MPORT_1_en_pipe_0;
  reg [3:0] mem_96_MPORT_1_addr_pipe_0;
  reg [7:0] mem_97 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_97_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_97_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_97_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_97_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_97_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_97_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_97_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_97_MPORT_1_en_pipe_0;
  reg [3:0] mem_97_MPORT_1_addr_pipe_0;
  reg [7:0] mem_98 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_98_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_98_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_98_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_98_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_98_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_98_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_98_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_98_MPORT_1_en_pipe_0;
  reg [3:0] mem_98_MPORT_1_addr_pipe_0;
  reg [7:0] mem_99 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_99_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_99_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_99_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_99_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_99_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_99_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_99_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_99_MPORT_1_en_pipe_0;
  reg [3:0] mem_99_MPORT_1_addr_pipe_0;
  reg [7:0] mem_100 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_100_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_100_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_100_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_100_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_100_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_100_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_100_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_100_MPORT_1_en_pipe_0;
  reg [3:0] mem_100_MPORT_1_addr_pipe_0;
  reg [7:0] mem_101 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_101_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_101_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_101_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_101_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_101_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_101_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_101_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_101_MPORT_1_en_pipe_0;
  reg [3:0] mem_101_MPORT_1_addr_pipe_0;
  reg [7:0] mem_102 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_102_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_102_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_102_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_102_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_102_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_102_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_102_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_102_MPORT_1_en_pipe_0;
  reg [3:0] mem_102_MPORT_1_addr_pipe_0;
  reg [7:0] mem_103 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_103_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_103_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_103_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_103_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_103_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_103_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_103_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_103_MPORT_1_en_pipe_0;
  reg [3:0] mem_103_MPORT_1_addr_pipe_0;
  reg [7:0] mem_104 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_104_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_104_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_104_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_104_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_104_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_104_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_104_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_104_MPORT_1_en_pipe_0;
  reg [3:0] mem_104_MPORT_1_addr_pipe_0;
  reg [7:0] mem_105 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_105_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_105_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_105_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_105_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_105_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_105_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_105_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_105_MPORT_1_en_pipe_0;
  reg [3:0] mem_105_MPORT_1_addr_pipe_0;
  reg [7:0] mem_106 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_106_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_106_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_106_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_106_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_106_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_106_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_106_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_106_MPORT_1_en_pipe_0;
  reg [3:0] mem_106_MPORT_1_addr_pipe_0;
  reg [7:0] mem_107 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_107_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_107_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_107_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_107_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_107_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_107_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_107_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_107_MPORT_1_en_pipe_0;
  reg [3:0] mem_107_MPORT_1_addr_pipe_0;
  reg [7:0] mem_108 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_108_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_108_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_108_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_108_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_108_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_108_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_108_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_108_MPORT_1_en_pipe_0;
  reg [3:0] mem_108_MPORT_1_addr_pipe_0;
  reg [7:0] mem_109 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_109_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_109_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_109_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_109_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_109_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_109_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_109_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_109_MPORT_1_en_pipe_0;
  reg [3:0] mem_109_MPORT_1_addr_pipe_0;
  reg [7:0] mem_110 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_110_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_110_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_110_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_110_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_110_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_110_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_110_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_110_MPORT_1_en_pipe_0;
  reg [3:0] mem_110_MPORT_1_addr_pipe_0;
  reg [7:0] mem_111 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_111_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_111_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_111_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_111_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_111_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_111_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_111_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_111_MPORT_1_en_pipe_0;
  reg [3:0] mem_111_MPORT_1_addr_pipe_0;
  reg [7:0] mem_112 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_112_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_112_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_112_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_112_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_112_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_112_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_112_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_112_MPORT_1_en_pipe_0;
  reg [3:0] mem_112_MPORT_1_addr_pipe_0;
  reg [7:0] mem_113 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_113_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_113_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_113_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_113_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_113_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_113_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_113_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_113_MPORT_1_en_pipe_0;
  reg [3:0] mem_113_MPORT_1_addr_pipe_0;
  reg [7:0] mem_114 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_114_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_114_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_114_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_114_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_114_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_114_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_114_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_114_MPORT_1_en_pipe_0;
  reg [3:0] mem_114_MPORT_1_addr_pipe_0;
  reg [7:0] mem_115 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_115_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_115_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_115_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_115_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_115_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_115_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_115_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_115_MPORT_1_en_pipe_0;
  reg [3:0] mem_115_MPORT_1_addr_pipe_0;
  reg [7:0] mem_116 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_116_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_116_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_116_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_116_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_116_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_116_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_116_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_116_MPORT_1_en_pipe_0;
  reg [3:0] mem_116_MPORT_1_addr_pipe_0;
  reg [7:0] mem_117 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_117_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_117_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_117_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_117_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_117_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_117_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_117_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_117_MPORT_1_en_pipe_0;
  reg [3:0] mem_117_MPORT_1_addr_pipe_0;
  reg [7:0] mem_118 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_118_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_118_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_118_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_118_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_118_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_118_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_118_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_118_MPORT_1_en_pipe_0;
  reg [3:0] mem_118_MPORT_1_addr_pipe_0;
  reg [7:0] mem_119 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_119_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_119_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_119_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_119_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_119_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_119_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_119_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_119_MPORT_1_en_pipe_0;
  reg [3:0] mem_119_MPORT_1_addr_pipe_0;
  reg [7:0] mem_120 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_120_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_120_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_120_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_120_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_120_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_120_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_120_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_120_MPORT_1_en_pipe_0;
  reg [3:0] mem_120_MPORT_1_addr_pipe_0;
  reg [7:0] mem_121 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_121_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_121_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_121_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_121_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_121_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_121_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_121_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_121_MPORT_1_en_pipe_0;
  reg [3:0] mem_121_MPORT_1_addr_pipe_0;
  reg [7:0] mem_122 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_122_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_122_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_122_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_122_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_122_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_122_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_122_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_122_MPORT_1_en_pipe_0;
  reg [3:0] mem_122_MPORT_1_addr_pipe_0;
  reg [7:0] mem_123 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_123_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_123_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_123_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_123_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_123_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_123_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_123_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_123_MPORT_1_en_pipe_0;
  reg [3:0] mem_123_MPORT_1_addr_pipe_0;
  reg [7:0] mem_124 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_124_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_124_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_124_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_124_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_124_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_124_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_124_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_124_MPORT_1_en_pipe_0;
  reg [3:0] mem_124_MPORT_1_addr_pipe_0;
  reg [7:0] mem_125 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_125_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_125_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_125_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_125_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_125_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_125_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_125_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_125_MPORT_1_en_pipe_0;
  reg [3:0] mem_125_MPORT_1_addr_pipe_0;
  reg [7:0] mem_126 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_126_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_126_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_126_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_126_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_126_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_126_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_126_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_126_MPORT_1_en_pipe_0;
  reg [3:0] mem_126_MPORT_1_addr_pipe_0;
  reg [7:0] mem_127 [0:15]; // @[BufferMemorySystem.scala 16:24]
  wire  mem_127_MPORT_1_en; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_127_MPORT_1_addr; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_127_MPORT_1_data; // @[BufferMemorySystem.scala 16:24]
  wire [7:0] mem_127_MPORT_data; // @[BufferMemorySystem.scala 16:24]
  wire [3:0] mem_127_MPORT_addr; // @[BufferMemorySystem.scala 16:24]
  wire  mem_127_MPORT_mask; // @[BufferMemorySystem.scala 16:24]
  wire  mem_127_MPORT_en; // @[BufferMemorySystem.scala 16:24]
  reg  mem_127_MPORT_1_en_pipe_0;
  reg [3:0] mem_127_MPORT_1_addr_pipe_0;
  reg [3:0] counter; // @[BufferMemorySystem.scala 14:24]
  wire [3:0] _counter_T_1 = counter + 4'h1; // @[BufferMemorySystem.scala 19:24]
  assign mem_0_MPORT_1_en = mem_0_MPORT_1_en_pipe_0;
  assign mem_0_MPORT_1_addr = mem_0_MPORT_1_addr_pipe_0;
  assign mem_0_MPORT_1_data = mem_0[mem_0_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_0_MPORT_data = io_adcValues_0;
  assign mem_0_MPORT_addr = counter;
  assign mem_0_MPORT_mask = 1'h1;
  assign mem_0_MPORT_en = 1'h1;
  assign mem_1_MPORT_1_en = mem_1_MPORT_1_en_pipe_0;
  assign mem_1_MPORT_1_addr = mem_1_MPORT_1_addr_pipe_0;
  assign mem_1_MPORT_1_data = mem_1[mem_1_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_1_MPORT_data = io_adcValues_1;
  assign mem_1_MPORT_addr = counter;
  assign mem_1_MPORT_mask = 1'h1;
  assign mem_1_MPORT_en = 1'h1;
  assign mem_2_MPORT_1_en = mem_2_MPORT_1_en_pipe_0;
  assign mem_2_MPORT_1_addr = mem_2_MPORT_1_addr_pipe_0;
  assign mem_2_MPORT_1_data = mem_2[mem_2_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_2_MPORT_data = io_adcValues_2;
  assign mem_2_MPORT_addr = counter;
  assign mem_2_MPORT_mask = 1'h1;
  assign mem_2_MPORT_en = 1'h1;
  assign mem_3_MPORT_1_en = mem_3_MPORT_1_en_pipe_0;
  assign mem_3_MPORT_1_addr = mem_3_MPORT_1_addr_pipe_0;
  assign mem_3_MPORT_1_data = mem_3[mem_3_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_3_MPORT_data = io_adcValues_3;
  assign mem_3_MPORT_addr = counter;
  assign mem_3_MPORT_mask = 1'h1;
  assign mem_3_MPORT_en = 1'h1;
  assign mem_4_MPORT_1_en = mem_4_MPORT_1_en_pipe_0;
  assign mem_4_MPORT_1_addr = mem_4_MPORT_1_addr_pipe_0;
  assign mem_4_MPORT_1_data = mem_4[mem_4_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_4_MPORT_data = io_adcValues_4;
  assign mem_4_MPORT_addr = counter;
  assign mem_4_MPORT_mask = 1'h1;
  assign mem_4_MPORT_en = 1'h1;
  assign mem_5_MPORT_1_en = mem_5_MPORT_1_en_pipe_0;
  assign mem_5_MPORT_1_addr = mem_5_MPORT_1_addr_pipe_0;
  assign mem_5_MPORT_1_data = mem_5[mem_5_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_5_MPORT_data = io_adcValues_5;
  assign mem_5_MPORT_addr = counter;
  assign mem_5_MPORT_mask = 1'h1;
  assign mem_5_MPORT_en = 1'h1;
  assign mem_6_MPORT_1_en = mem_6_MPORT_1_en_pipe_0;
  assign mem_6_MPORT_1_addr = mem_6_MPORT_1_addr_pipe_0;
  assign mem_6_MPORT_1_data = mem_6[mem_6_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_6_MPORT_data = io_adcValues_6;
  assign mem_6_MPORT_addr = counter;
  assign mem_6_MPORT_mask = 1'h1;
  assign mem_6_MPORT_en = 1'h1;
  assign mem_7_MPORT_1_en = mem_7_MPORT_1_en_pipe_0;
  assign mem_7_MPORT_1_addr = mem_7_MPORT_1_addr_pipe_0;
  assign mem_7_MPORT_1_data = mem_7[mem_7_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_7_MPORT_data = io_adcValues_7;
  assign mem_7_MPORT_addr = counter;
  assign mem_7_MPORT_mask = 1'h1;
  assign mem_7_MPORT_en = 1'h1;
  assign mem_8_MPORT_1_en = mem_8_MPORT_1_en_pipe_0;
  assign mem_8_MPORT_1_addr = mem_8_MPORT_1_addr_pipe_0;
  assign mem_8_MPORT_1_data = mem_8[mem_8_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_8_MPORT_data = io_adcValues_8;
  assign mem_8_MPORT_addr = counter;
  assign mem_8_MPORT_mask = 1'h1;
  assign mem_8_MPORT_en = 1'h1;
  assign mem_9_MPORT_1_en = mem_9_MPORT_1_en_pipe_0;
  assign mem_9_MPORT_1_addr = mem_9_MPORT_1_addr_pipe_0;
  assign mem_9_MPORT_1_data = mem_9[mem_9_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_9_MPORT_data = io_adcValues_9;
  assign mem_9_MPORT_addr = counter;
  assign mem_9_MPORT_mask = 1'h1;
  assign mem_9_MPORT_en = 1'h1;
  assign mem_10_MPORT_1_en = mem_10_MPORT_1_en_pipe_0;
  assign mem_10_MPORT_1_addr = mem_10_MPORT_1_addr_pipe_0;
  assign mem_10_MPORT_1_data = mem_10[mem_10_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_10_MPORT_data = io_adcValues_10;
  assign mem_10_MPORT_addr = counter;
  assign mem_10_MPORT_mask = 1'h1;
  assign mem_10_MPORT_en = 1'h1;
  assign mem_11_MPORT_1_en = mem_11_MPORT_1_en_pipe_0;
  assign mem_11_MPORT_1_addr = mem_11_MPORT_1_addr_pipe_0;
  assign mem_11_MPORT_1_data = mem_11[mem_11_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_11_MPORT_data = io_adcValues_11;
  assign mem_11_MPORT_addr = counter;
  assign mem_11_MPORT_mask = 1'h1;
  assign mem_11_MPORT_en = 1'h1;
  assign mem_12_MPORT_1_en = mem_12_MPORT_1_en_pipe_0;
  assign mem_12_MPORT_1_addr = mem_12_MPORT_1_addr_pipe_0;
  assign mem_12_MPORT_1_data = mem_12[mem_12_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_12_MPORT_data = io_adcValues_12;
  assign mem_12_MPORT_addr = counter;
  assign mem_12_MPORT_mask = 1'h1;
  assign mem_12_MPORT_en = 1'h1;
  assign mem_13_MPORT_1_en = mem_13_MPORT_1_en_pipe_0;
  assign mem_13_MPORT_1_addr = mem_13_MPORT_1_addr_pipe_0;
  assign mem_13_MPORT_1_data = mem_13[mem_13_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_13_MPORT_data = io_adcValues_13;
  assign mem_13_MPORT_addr = counter;
  assign mem_13_MPORT_mask = 1'h1;
  assign mem_13_MPORT_en = 1'h1;
  assign mem_14_MPORT_1_en = mem_14_MPORT_1_en_pipe_0;
  assign mem_14_MPORT_1_addr = mem_14_MPORT_1_addr_pipe_0;
  assign mem_14_MPORT_1_data = mem_14[mem_14_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_14_MPORT_data = io_adcValues_14;
  assign mem_14_MPORT_addr = counter;
  assign mem_14_MPORT_mask = 1'h1;
  assign mem_14_MPORT_en = 1'h1;
  assign mem_15_MPORT_1_en = mem_15_MPORT_1_en_pipe_0;
  assign mem_15_MPORT_1_addr = mem_15_MPORT_1_addr_pipe_0;
  assign mem_15_MPORT_1_data = mem_15[mem_15_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_15_MPORT_data = io_adcValues_15;
  assign mem_15_MPORT_addr = counter;
  assign mem_15_MPORT_mask = 1'h1;
  assign mem_15_MPORT_en = 1'h1;
  assign mem_16_MPORT_1_en = mem_16_MPORT_1_en_pipe_0;
  assign mem_16_MPORT_1_addr = mem_16_MPORT_1_addr_pipe_0;
  assign mem_16_MPORT_1_data = mem_16[mem_16_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_16_MPORT_data = io_adcValues_16;
  assign mem_16_MPORT_addr = counter;
  assign mem_16_MPORT_mask = 1'h1;
  assign mem_16_MPORT_en = 1'h1;
  assign mem_17_MPORT_1_en = mem_17_MPORT_1_en_pipe_0;
  assign mem_17_MPORT_1_addr = mem_17_MPORT_1_addr_pipe_0;
  assign mem_17_MPORT_1_data = mem_17[mem_17_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_17_MPORT_data = io_adcValues_17;
  assign mem_17_MPORT_addr = counter;
  assign mem_17_MPORT_mask = 1'h1;
  assign mem_17_MPORT_en = 1'h1;
  assign mem_18_MPORT_1_en = mem_18_MPORT_1_en_pipe_0;
  assign mem_18_MPORT_1_addr = mem_18_MPORT_1_addr_pipe_0;
  assign mem_18_MPORT_1_data = mem_18[mem_18_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_18_MPORT_data = io_adcValues_18;
  assign mem_18_MPORT_addr = counter;
  assign mem_18_MPORT_mask = 1'h1;
  assign mem_18_MPORT_en = 1'h1;
  assign mem_19_MPORT_1_en = mem_19_MPORT_1_en_pipe_0;
  assign mem_19_MPORT_1_addr = mem_19_MPORT_1_addr_pipe_0;
  assign mem_19_MPORT_1_data = mem_19[mem_19_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_19_MPORT_data = io_adcValues_19;
  assign mem_19_MPORT_addr = counter;
  assign mem_19_MPORT_mask = 1'h1;
  assign mem_19_MPORT_en = 1'h1;
  assign mem_20_MPORT_1_en = mem_20_MPORT_1_en_pipe_0;
  assign mem_20_MPORT_1_addr = mem_20_MPORT_1_addr_pipe_0;
  assign mem_20_MPORT_1_data = mem_20[mem_20_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_20_MPORT_data = io_adcValues_20;
  assign mem_20_MPORT_addr = counter;
  assign mem_20_MPORT_mask = 1'h1;
  assign mem_20_MPORT_en = 1'h1;
  assign mem_21_MPORT_1_en = mem_21_MPORT_1_en_pipe_0;
  assign mem_21_MPORT_1_addr = mem_21_MPORT_1_addr_pipe_0;
  assign mem_21_MPORT_1_data = mem_21[mem_21_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_21_MPORT_data = io_adcValues_21;
  assign mem_21_MPORT_addr = counter;
  assign mem_21_MPORT_mask = 1'h1;
  assign mem_21_MPORT_en = 1'h1;
  assign mem_22_MPORT_1_en = mem_22_MPORT_1_en_pipe_0;
  assign mem_22_MPORT_1_addr = mem_22_MPORT_1_addr_pipe_0;
  assign mem_22_MPORT_1_data = mem_22[mem_22_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_22_MPORT_data = io_adcValues_22;
  assign mem_22_MPORT_addr = counter;
  assign mem_22_MPORT_mask = 1'h1;
  assign mem_22_MPORT_en = 1'h1;
  assign mem_23_MPORT_1_en = mem_23_MPORT_1_en_pipe_0;
  assign mem_23_MPORT_1_addr = mem_23_MPORT_1_addr_pipe_0;
  assign mem_23_MPORT_1_data = mem_23[mem_23_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_23_MPORT_data = io_adcValues_23;
  assign mem_23_MPORT_addr = counter;
  assign mem_23_MPORT_mask = 1'h1;
  assign mem_23_MPORT_en = 1'h1;
  assign mem_24_MPORT_1_en = mem_24_MPORT_1_en_pipe_0;
  assign mem_24_MPORT_1_addr = mem_24_MPORT_1_addr_pipe_0;
  assign mem_24_MPORT_1_data = mem_24[mem_24_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_24_MPORT_data = io_adcValues_24;
  assign mem_24_MPORT_addr = counter;
  assign mem_24_MPORT_mask = 1'h1;
  assign mem_24_MPORT_en = 1'h1;
  assign mem_25_MPORT_1_en = mem_25_MPORT_1_en_pipe_0;
  assign mem_25_MPORT_1_addr = mem_25_MPORT_1_addr_pipe_0;
  assign mem_25_MPORT_1_data = mem_25[mem_25_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_25_MPORT_data = io_adcValues_25;
  assign mem_25_MPORT_addr = counter;
  assign mem_25_MPORT_mask = 1'h1;
  assign mem_25_MPORT_en = 1'h1;
  assign mem_26_MPORT_1_en = mem_26_MPORT_1_en_pipe_0;
  assign mem_26_MPORT_1_addr = mem_26_MPORT_1_addr_pipe_0;
  assign mem_26_MPORT_1_data = mem_26[mem_26_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_26_MPORT_data = io_adcValues_26;
  assign mem_26_MPORT_addr = counter;
  assign mem_26_MPORT_mask = 1'h1;
  assign mem_26_MPORT_en = 1'h1;
  assign mem_27_MPORT_1_en = mem_27_MPORT_1_en_pipe_0;
  assign mem_27_MPORT_1_addr = mem_27_MPORT_1_addr_pipe_0;
  assign mem_27_MPORT_1_data = mem_27[mem_27_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_27_MPORT_data = io_adcValues_27;
  assign mem_27_MPORT_addr = counter;
  assign mem_27_MPORT_mask = 1'h1;
  assign mem_27_MPORT_en = 1'h1;
  assign mem_28_MPORT_1_en = mem_28_MPORT_1_en_pipe_0;
  assign mem_28_MPORT_1_addr = mem_28_MPORT_1_addr_pipe_0;
  assign mem_28_MPORT_1_data = mem_28[mem_28_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_28_MPORT_data = io_adcValues_28;
  assign mem_28_MPORT_addr = counter;
  assign mem_28_MPORT_mask = 1'h1;
  assign mem_28_MPORT_en = 1'h1;
  assign mem_29_MPORT_1_en = mem_29_MPORT_1_en_pipe_0;
  assign mem_29_MPORT_1_addr = mem_29_MPORT_1_addr_pipe_0;
  assign mem_29_MPORT_1_data = mem_29[mem_29_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_29_MPORT_data = io_adcValues_29;
  assign mem_29_MPORT_addr = counter;
  assign mem_29_MPORT_mask = 1'h1;
  assign mem_29_MPORT_en = 1'h1;
  assign mem_30_MPORT_1_en = mem_30_MPORT_1_en_pipe_0;
  assign mem_30_MPORT_1_addr = mem_30_MPORT_1_addr_pipe_0;
  assign mem_30_MPORT_1_data = mem_30[mem_30_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_30_MPORT_data = io_adcValues_30;
  assign mem_30_MPORT_addr = counter;
  assign mem_30_MPORT_mask = 1'h1;
  assign mem_30_MPORT_en = 1'h1;
  assign mem_31_MPORT_1_en = mem_31_MPORT_1_en_pipe_0;
  assign mem_31_MPORT_1_addr = mem_31_MPORT_1_addr_pipe_0;
  assign mem_31_MPORT_1_data = mem_31[mem_31_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_31_MPORT_data = io_adcValues_31;
  assign mem_31_MPORT_addr = counter;
  assign mem_31_MPORT_mask = 1'h1;
  assign mem_31_MPORT_en = 1'h1;
  assign mem_32_MPORT_1_en = mem_32_MPORT_1_en_pipe_0;
  assign mem_32_MPORT_1_addr = mem_32_MPORT_1_addr_pipe_0;
  assign mem_32_MPORT_1_data = mem_32[mem_32_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_32_MPORT_data = io_adcValues_32;
  assign mem_32_MPORT_addr = counter;
  assign mem_32_MPORT_mask = 1'h1;
  assign mem_32_MPORT_en = 1'h1;
  assign mem_33_MPORT_1_en = mem_33_MPORT_1_en_pipe_0;
  assign mem_33_MPORT_1_addr = mem_33_MPORT_1_addr_pipe_0;
  assign mem_33_MPORT_1_data = mem_33[mem_33_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_33_MPORT_data = io_adcValues_33;
  assign mem_33_MPORT_addr = counter;
  assign mem_33_MPORT_mask = 1'h1;
  assign mem_33_MPORT_en = 1'h1;
  assign mem_34_MPORT_1_en = mem_34_MPORT_1_en_pipe_0;
  assign mem_34_MPORT_1_addr = mem_34_MPORT_1_addr_pipe_0;
  assign mem_34_MPORT_1_data = mem_34[mem_34_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_34_MPORT_data = io_adcValues_34;
  assign mem_34_MPORT_addr = counter;
  assign mem_34_MPORT_mask = 1'h1;
  assign mem_34_MPORT_en = 1'h1;
  assign mem_35_MPORT_1_en = mem_35_MPORT_1_en_pipe_0;
  assign mem_35_MPORT_1_addr = mem_35_MPORT_1_addr_pipe_0;
  assign mem_35_MPORT_1_data = mem_35[mem_35_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_35_MPORT_data = io_adcValues_35;
  assign mem_35_MPORT_addr = counter;
  assign mem_35_MPORT_mask = 1'h1;
  assign mem_35_MPORT_en = 1'h1;
  assign mem_36_MPORT_1_en = mem_36_MPORT_1_en_pipe_0;
  assign mem_36_MPORT_1_addr = mem_36_MPORT_1_addr_pipe_0;
  assign mem_36_MPORT_1_data = mem_36[mem_36_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_36_MPORT_data = io_adcValues_36;
  assign mem_36_MPORT_addr = counter;
  assign mem_36_MPORT_mask = 1'h1;
  assign mem_36_MPORT_en = 1'h1;
  assign mem_37_MPORT_1_en = mem_37_MPORT_1_en_pipe_0;
  assign mem_37_MPORT_1_addr = mem_37_MPORT_1_addr_pipe_0;
  assign mem_37_MPORT_1_data = mem_37[mem_37_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_37_MPORT_data = io_adcValues_37;
  assign mem_37_MPORT_addr = counter;
  assign mem_37_MPORT_mask = 1'h1;
  assign mem_37_MPORT_en = 1'h1;
  assign mem_38_MPORT_1_en = mem_38_MPORT_1_en_pipe_0;
  assign mem_38_MPORT_1_addr = mem_38_MPORT_1_addr_pipe_0;
  assign mem_38_MPORT_1_data = mem_38[mem_38_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_38_MPORT_data = io_adcValues_38;
  assign mem_38_MPORT_addr = counter;
  assign mem_38_MPORT_mask = 1'h1;
  assign mem_38_MPORT_en = 1'h1;
  assign mem_39_MPORT_1_en = mem_39_MPORT_1_en_pipe_0;
  assign mem_39_MPORT_1_addr = mem_39_MPORT_1_addr_pipe_0;
  assign mem_39_MPORT_1_data = mem_39[mem_39_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_39_MPORT_data = io_adcValues_39;
  assign mem_39_MPORT_addr = counter;
  assign mem_39_MPORT_mask = 1'h1;
  assign mem_39_MPORT_en = 1'h1;
  assign mem_40_MPORT_1_en = mem_40_MPORT_1_en_pipe_0;
  assign mem_40_MPORT_1_addr = mem_40_MPORT_1_addr_pipe_0;
  assign mem_40_MPORT_1_data = mem_40[mem_40_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_40_MPORT_data = io_adcValues_40;
  assign mem_40_MPORT_addr = counter;
  assign mem_40_MPORT_mask = 1'h1;
  assign mem_40_MPORT_en = 1'h1;
  assign mem_41_MPORT_1_en = mem_41_MPORT_1_en_pipe_0;
  assign mem_41_MPORT_1_addr = mem_41_MPORT_1_addr_pipe_0;
  assign mem_41_MPORT_1_data = mem_41[mem_41_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_41_MPORT_data = io_adcValues_41;
  assign mem_41_MPORT_addr = counter;
  assign mem_41_MPORT_mask = 1'h1;
  assign mem_41_MPORT_en = 1'h1;
  assign mem_42_MPORT_1_en = mem_42_MPORT_1_en_pipe_0;
  assign mem_42_MPORT_1_addr = mem_42_MPORT_1_addr_pipe_0;
  assign mem_42_MPORT_1_data = mem_42[mem_42_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_42_MPORT_data = io_adcValues_42;
  assign mem_42_MPORT_addr = counter;
  assign mem_42_MPORT_mask = 1'h1;
  assign mem_42_MPORT_en = 1'h1;
  assign mem_43_MPORT_1_en = mem_43_MPORT_1_en_pipe_0;
  assign mem_43_MPORT_1_addr = mem_43_MPORT_1_addr_pipe_0;
  assign mem_43_MPORT_1_data = mem_43[mem_43_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_43_MPORT_data = io_adcValues_43;
  assign mem_43_MPORT_addr = counter;
  assign mem_43_MPORT_mask = 1'h1;
  assign mem_43_MPORT_en = 1'h1;
  assign mem_44_MPORT_1_en = mem_44_MPORT_1_en_pipe_0;
  assign mem_44_MPORT_1_addr = mem_44_MPORT_1_addr_pipe_0;
  assign mem_44_MPORT_1_data = mem_44[mem_44_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_44_MPORT_data = io_adcValues_44;
  assign mem_44_MPORT_addr = counter;
  assign mem_44_MPORT_mask = 1'h1;
  assign mem_44_MPORT_en = 1'h1;
  assign mem_45_MPORT_1_en = mem_45_MPORT_1_en_pipe_0;
  assign mem_45_MPORT_1_addr = mem_45_MPORT_1_addr_pipe_0;
  assign mem_45_MPORT_1_data = mem_45[mem_45_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_45_MPORT_data = io_adcValues_45;
  assign mem_45_MPORT_addr = counter;
  assign mem_45_MPORT_mask = 1'h1;
  assign mem_45_MPORT_en = 1'h1;
  assign mem_46_MPORT_1_en = mem_46_MPORT_1_en_pipe_0;
  assign mem_46_MPORT_1_addr = mem_46_MPORT_1_addr_pipe_0;
  assign mem_46_MPORT_1_data = mem_46[mem_46_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_46_MPORT_data = io_adcValues_46;
  assign mem_46_MPORT_addr = counter;
  assign mem_46_MPORT_mask = 1'h1;
  assign mem_46_MPORT_en = 1'h1;
  assign mem_47_MPORT_1_en = mem_47_MPORT_1_en_pipe_0;
  assign mem_47_MPORT_1_addr = mem_47_MPORT_1_addr_pipe_0;
  assign mem_47_MPORT_1_data = mem_47[mem_47_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_47_MPORT_data = io_adcValues_47;
  assign mem_47_MPORT_addr = counter;
  assign mem_47_MPORT_mask = 1'h1;
  assign mem_47_MPORT_en = 1'h1;
  assign mem_48_MPORT_1_en = mem_48_MPORT_1_en_pipe_0;
  assign mem_48_MPORT_1_addr = mem_48_MPORT_1_addr_pipe_0;
  assign mem_48_MPORT_1_data = mem_48[mem_48_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_48_MPORT_data = io_adcValues_48;
  assign mem_48_MPORT_addr = counter;
  assign mem_48_MPORT_mask = 1'h1;
  assign mem_48_MPORT_en = 1'h1;
  assign mem_49_MPORT_1_en = mem_49_MPORT_1_en_pipe_0;
  assign mem_49_MPORT_1_addr = mem_49_MPORT_1_addr_pipe_0;
  assign mem_49_MPORT_1_data = mem_49[mem_49_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_49_MPORT_data = io_adcValues_49;
  assign mem_49_MPORT_addr = counter;
  assign mem_49_MPORT_mask = 1'h1;
  assign mem_49_MPORT_en = 1'h1;
  assign mem_50_MPORT_1_en = mem_50_MPORT_1_en_pipe_0;
  assign mem_50_MPORT_1_addr = mem_50_MPORT_1_addr_pipe_0;
  assign mem_50_MPORT_1_data = mem_50[mem_50_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_50_MPORT_data = io_adcValues_50;
  assign mem_50_MPORT_addr = counter;
  assign mem_50_MPORT_mask = 1'h1;
  assign mem_50_MPORT_en = 1'h1;
  assign mem_51_MPORT_1_en = mem_51_MPORT_1_en_pipe_0;
  assign mem_51_MPORT_1_addr = mem_51_MPORT_1_addr_pipe_0;
  assign mem_51_MPORT_1_data = mem_51[mem_51_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_51_MPORT_data = io_adcValues_51;
  assign mem_51_MPORT_addr = counter;
  assign mem_51_MPORT_mask = 1'h1;
  assign mem_51_MPORT_en = 1'h1;
  assign mem_52_MPORT_1_en = mem_52_MPORT_1_en_pipe_0;
  assign mem_52_MPORT_1_addr = mem_52_MPORT_1_addr_pipe_0;
  assign mem_52_MPORT_1_data = mem_52[mem_52_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_52_MPORT_data = io_adcValues_52;
  assign mem_52_MPORT_addr = counter;
  assign mem_52_MPORT_mask = 1'h1;
  assign mem_52_MPORT_en = 1'h1;
  assign mem_53_MPORT_1_en = mem_53_MPORT_1_en_pipe_0;
  assign mem_53_MPORT_1_addr = mem_53_MPORT_1_addr_pipe_0;
  assign mem_53_MPORT_1_data = mem_53[mem_53_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_53_MPORT_data = io_adcValues_53;
  assign mem_53_MPORT_addr = counter;
  assign mem_53_MPORT_mask = 1'h1;
  assign mem_53_MPORT_en = 1'h1;
  assign mem_54_MPORT_1_en = mem_54_MPORT_1_en_pipe_0;
  assign mem_54_MPORT_1_addr = mem_54_MPORT_1_addr_pipe_0;
  assign mem_54_MPORT_1_data = mem_54[mem_54_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_54_MPORT_data = io_adcValues_54;
  assign mem_54_MPORT_addr = counter;
  assign mem_54_MPORT_mask = 1'h1;
  assign mem_54_MPORT_en = 1'h1;
  assign mem_55_MPORT_1_en = mem_55_MPORT_1_en_pipe_0;
  assign mem_55_MPORT_1_addr = mem_55_MPORT_1_addr_pipe_0;
  assign mem_55_MPORT_1_data = mem_55[mem_55_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_55_MPORT_data = io_adcValues_55;
  assign mem_55_MPORT_addr = counter;
  assign mem_55_MPORT_mask = 1'h1;
  assign mem_55_MPORT_en = 1'h1;
  assign mem_56_MPORT_1_en = mem_56_MPORT_1_en_pipe_0;
  assign mem_56_MPORT_1_addr = mem_56_MPORT_1_addr_pipe_0;
  assign mem_56_MPORT_1_data = mem_56[mem_56_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_56_MPORT_data = io_adcValues_56;
  assign mem_56_MPORT_addr = counter;
  assign mem_56_MPORT_mask = 1'h1;
  assign mem_56_MPORT_en = 1'h1;
  assign mem_57_MPORT_1_en = mem_57_MPORT_1_en_pipe_0;
  assign mem_57_MPORT_1_addr = mem_57_MPORT_1_addr_pipe_0;
  assign mem_57_MPORT_1_data = mem_57[mem_57_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_57_MPORT_data = io_adcValues_57;
  assign mem_57_MPORT_addr = counter;
  assign mem_57_MPORT_mask = 1'h1;
  assign mem_57_MPORT_en = 1'h1;
  assign mem_58_MPORT_1_en = mem_58_MPORT_1_en_pipe_0;
  assign mem_58_MPORT_1_addr = mem_58_MPORT_1_addr_pipe_0;
  assign mem_58_MPORT_1_data = mem_58[mem_58_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_58_MPORT_data = io_adcValues_58;
  assign mem_58_MPORT_addr = counter;
  assign mem_58_MPORT_mask = 1'h1;
  assign mem_58_MPORT_en = 1'h1;
  assign mem_59_MPORT_1_en = mem_59_MPORT_1_en_pipe_0;
  assign mem_59_MPORT_1_addr = mem_59_MPORT_1_addr_pipe_0;
  assign mem_59_MPORT_1_data = mem_59[mem_59_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_59_MPORT_data = io_adcValues_59;
  assign mem_59_MPORT_addr = counter;
  assign mem_59_MPORT_mask = 1'h1;
  assign mem_59_MPORT_en = 1'h1;
  assign mem_60_MPORT_1_en = mem_60_MPORT_1_en_pipe_0;
  assign mem_60_MPORT_1_addr = mem_60_MPORT_1_addr_pipe_0;
  assign mem_60_MPORT_1_data = mem_60[mem_60_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_60_MPORT_data = io_adcValues_60;
  assign mem_60_MPORT_addr = counter;
  assign mem_60_MPORT_mask = 1'h1;
  assign mem_60_MPORT_en = 1'h1;
  assign mem_61_MPORT_1_en = mem_61_MPORT_1_en_pipe_0;
  assign mem_61_MPORT_1_addr = mem_61_MPORT_1_addr_pipe_0;
  assign mem_61_MPORT_1_data = mem_61[mem_61_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_61_MPORT_data = io_adcValues_61;
  assign mem_61_MPORT_addr = counter;
  assign mem_61_MPORT_mask = 1'h1;
  assign mem_61_MPORT_en = 1'h1;
  assign mem_62_MPORT_1_en = mem_62_MPORT_1_en_pipe_0;
  assign mem_62_MPORT_1_addr = mem_62_MPORT_1_addr_pipe_0;
  assign mem_62_MPORT_1_data = mem_62[mem_62_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_62_MPORT_data = io_adcValues_62;
  assign mem_62_MPORT_addr = counter;
  assign mem_62_MPORT_mask = 1'h1;
  assign mem_62_MPORT_en = 1'h1;
  assign mem_63_MPORT_1_en = mem_63_MPORT_1_en_pipe_0;
  assign mem_63_MPORT_1_addr = mem_63_MPORT_1_addr_pipe_0;
  assign mem_63_MPORT_1_data = mem_63[mem_63_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_63_MPORT_data = io_adcValues_63;
  assign mem_63_MPORT_addr = counter;
  assign mem_63_MPORT_mask = 1'h1;
  assign mem_63_MPORT_en = 1'h1;
  assign mem_64_MPORT_1_en = mem_64_MPORT_1_en_pipe_0;
  assign mem_64_MPORT_1_addr = mem_64_MPORT_1_addr_pipe_0;
  assign mem_64_MPORT_1_data = mem_64[mem_64_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_64_MPORT_data = io_adcValues_64;
  assign mem_64_MPORT_addr = counter;
  assign mem_64_MPORT_mask = 1'h1;
  assign mem_64_MPORT_en = 1'h1;
  assign mem_65_MPORT_1_en = mem_65_MPORT_1_en_pipe_0;
  assign mem_65_MPORT_1_addr = mem_65_MPORT_1_addr_pipe_0;
  assign mem_65_MPORT_1_data = mem_65[mem_65_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_65_MPORT_data = io_adcValues_65;
  assign mem_65_MPORT_addr = counter;
  assign mem_65_MPORT_mask = 1'h1;
  assign mem_65_MPORT_en = 1'h1;
  assign mem_66_MPORT_1_en = mem_66_MPORT_1_en_pipe_0;
  assign mem_66_MPORT_1_addr = mem_66_MPORT_1_addr_pipe_0;
  assign mem_66_MPORT_1_data = mem_66[mem_66_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_66_MPORT_data = io_adcValues_66;
  assign mem_66_MPORT_addr = counter;
  assign mem_66_MPORT_mask = 1'h1;
  assign mem_66_MPORT_en = 1'h1;
  assign mem_67_MPORT_1_en = mem_67_MPORT_1_en_pipe_0;
  assign mem_67_MPORT_1_addr = mem_67_MPORT_1_addr_pipe_0;
  assign mem_67_MPORT_1_data = mem_67[mem_67_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_67_MPORT_data = io_adcValues_67;
  assign mem_67_MPORT_addr = counter;
  assign mem_67_MPORT_mask = 1'h1;
  assign mem_67_MPORT_en = 1'h1;
  assign mem_68_MPORT_1_en = mem_68_MPORT_1_en_pipe_0;
  assign mem_68_MPORT_1_addr = mem_68_MPORT_1_addr_pipe_0;
  assign mem_68_MPORT_1_data = mem_68[mem_68_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_68_MPORT_data = io_adcValues_68;
  assign mem_68_MPORT_addr = counter;
  assign mem_68_MPORT_mask = 1'h1;
  assign mem_68_MPORT_en = 1'h1;
  assign mem_69_MPORT_1_en = mem_69_MPORT_1_en_pipe_0;
  assign mem_69_MPORT_1_addr = mem_69_MPORT_1_addr_pipe_0;
  assign mem_69_MPORT_1_data = mem_69[mem_69_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_69_MPORT_data = io_adcValues_69;
  assign mem_69_MPORT_addr = counter;
  assign mem_69_MPORT_mask = 1'h1;
  assign mem_69_MPORT_en = 1'h1;
  assign mem_70_MPORT_1_en = mem_70_MPORT_1_en_pipe_0;
  assign mem_70_MPORT_1_addr = mem_70_MPORT_1_addr_pipe_0;
  assign mem_70_MPORT_1_data = mem_70[mem_70_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_70_MPORT_data = io_adcValues_70;
  assign mem_70_MPORT_addr = counter;
  assign mem_70_MPORT_mask = 1'h1;
  assign mem_70_MPORT_en = 1'h1;
  assign mem_71_MPORT_1_en = mem_71_MPORT_1_en_pipe_0;
  assign mem_71_MPORT_1_addr = mem_71_MPORT_1_addr_pipe_0;
  assign mem_71_MPORT_1_data = mem_71[mem_71_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_71_MPORT_data = io_adcValues_71;
  assign mem_71_MPORT_addr = counter;
  assign mem_71_MPORT_mask = 1'h1;
  assign mem_71_MPORT_en = 1'h1;
  assign mem_72_MPORT_1_en = mem_72_MPORT_1_en_pipe_0;
  assign mem_72_MPORT_1_addr = mem_72_MPORT_1_addr_pipe_0;
  assign mem_72_MPORT_1_data = mem_72[mem_72_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_72_MPORT_data = io_adcValues_72;
  assign mem_72_MPORT_addr = counter;
  assign mem_72_MPORT_mask = 1'h1;
  assign mem_72_MPORT_en = 1'h1;
  assign mem_73_MPORT_1_en = mem_73_MPORT_1_en_pipe_0;
  assign mem_73_MPORT_1_addr = mem_73_MPORT_1_addr_pipe_0;
  assign mem_73_MPORT_1_data = mem_73[mem_73_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_73_MPORT_data = io_adcValues_73;
  assign mem_73_MPORT_addr = counter;
  assign mem_73_MPORT_mask = 1'h1;
  assign mem_73_MPORT_en = 1'h1;
  assign mem_74_MPORT_1_en = mem_74_MPORT_1_en_pipe_0;
  assign mem_74_MPORT_1_addr = mem_74_MPORT_1_addr_pipe_0;
  assign mem_74_MPORT_1_data = mem_74[mem_74_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_74_MPORT_data = io_adcValues_74;
  assign mem_74_MPORT_addr = counter;
  assign mem_74_MPORT_mask = 1'h1;
  assign mem_74_MPORT_en = 1'h1;
  assign mem_75_MPORT_1_en = mem_75_MPORT_1_en_pipe_0;
  assign mem_75_MPORT_1_addr = mem_75_MPORT_1_addr_pipe_0;
  assign mem_75_MPORT_1_data = mem_75[mem_75_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_75_MPORT_data = io_adcValues_75;
  assign mem_75_MPORT_addr = counter;
  assign mem_75_MPORT_mask = 1'h1;
  assign mem_75_MPORT_en = 1'h1;
  assign mem_76_MPORT_1_en = mem_76_MPORT_1_en_pipe_0;
  assign mem_76_MPORT_1_addr = mem_76_MPORT_1_addr_pipe_0;
  assign mem_76_MPORT_1_data = mem_76[mem_76_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_76_MPORT_data = io_adcValues_76;
  assign mem_76_MPORT_addr = counter;
  assign mem_76_MPORT_mask = 1'h1;
  assign mem_76_MPORT_en = 1'h1;
  assign mem_77_MPORT_1_en = mem_77_MPORT_1_en_pipe_0;
  assign mem_77_MPORT_1_addr = mem_77_MPORT_1_addr_pipe_0;
  assign mem_77_MPORT_1_data = mem_77[mem_77_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_77_MPORT_data = io_adcValues_77;
  assign mem_77_MPORT_addr = counter;
  assign mem_77_MPORT_mask = 1'h1;
  assign mem_77_MPORT_en = 1'h1;
  assign mem_78_MPORT_1_en = mem_78_MPORT_1_en_pipe_0;
  assign mem_78_MPORT_1_addr = mem_78_MPORT_1_addr_pipe_0;
  assign mem_78_MPORT_1_data = mem_78[mem_78_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_78_MPORT_data = io_adcValues_78;
  assign mem_78_MPORT_addr = counter;
  assign mem_78_MPORT_mask = 1'h1;
  assign mem_78_MPORT_en = 1'h1;
  assign mem_79_MPORT_1_en = mem_79_MPORT_1_en_pipe_0;
  assign mem_79_MPORT_1_addr = mem_79_MPORT_1_addr_pipe_0;
  assign mem_79_MPORT_1_data = mem_79[mem_79_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_79_MPORT_data = io_adcValues_79;
  assign mem_79_MPORT_addr = counter;
  assign mem_79_MPORT_mask = 1'h1;
  assign mem_79_MPORT_en = 1'h1;
  assign mem_80_MPORT_1_en = mem_80_MPORT_1_en_pipe_0;
  assign mem_80_MPORT_1_addr = mem_80_MPORT_1_addr_pipe_0;
  assign mem_80_MPORT_1_data = mem_80[mem_80_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_80_MPORT_data = io_adcValues_80;
  assign mem_80_MPORT_addr = counter;
  assign mem_80_MPORT_mask = 1'h1;
  assign mem_80_MPORT_en = 1'h1;
  assign mem_81_MPORT_1_en = mem_81_MPORT_1_en_pipe_0;
  assign mem_81_MPORT_1_addr = mem_81_MPORT_1_addr_pipe_0;
  assign mem_81_MPORT_1_data = mem_81[mem_81_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_81_MPORT_data = io_adcValues_81;
  assign mem_81_MPORT_addr = counter;
  assign mem_81_MPORT_mask = 1'h1;
  assign mem_81_MPORT_en = 1'h1;
  assign mem_82_MPORT_1_en = mem_82_MPORT_1_en_pipe_0;
  assign mem_82_MPORT_1_addr = mem_82_MPORT_1_addr_pipe_0;
  assign mem_82_MPORT_1_data = mem_82[mem_82_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_82_MPORT_data = io_adcValues_82;
  assign mem_82_MPORT_addr = counter;
  assign mem_82_MPORT_mask = 1'h1;
  assign mem_82_MPORT_en = 1'h1;
  assign mem_83_MPORT_1_en = mem_83_MPORT_1_en_pipe_0;
  assign mem_83_MPORT_1_addr = mem_83_MPORT_1_addr_pipe_0;
  assign mem_83_MPORT_1_data = mem_83[mem_83_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_83_MPORT_data = io_adcValues_83;
  assign mem_83_MPORT_addr = counter;
  assign mem_83_MPORT_mask = 1'h1;
  assign mem_83_MPORT_en = 1'h1;
  assign mem_84_MPORT_1_en = mem_84_MPORT_1_en_pipe_0;
  assign mem_84_MPORT_1_addr = mem_84_MPORT_1_addr_pipe_0;
  assign mem_84_MPORT_1_data = mem_84[mem_84_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_84_MPORT_data = io_adcValues_84;
  assign mem_84_MPORT_addr = counter;
  assign mem_84_MPORT_mask = 1'h1;
  assign mem_84_MPORT_en = 1'h1;
  assign mem_85_MPORT_1_en = mem_85_MPORT_1_en_pipe_0;
  assign mem_85_MPORT_1_addr = mem_85_MPORT_1_addr_pipe_0;
  assign mem_85_MPORT_1_data = mem_85[mem_85_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_85_MPORT_data = io_adcValues_85;
  assign mem_85_MPORT_addr = counter;
  assign mem_85_MPORT_mask = 1'h1;
  assign mem_85_MPORT_en = 1'h1;
  assign mem_86_MPORT_1_en = mem_86_MPORT_1_en_pipe_0;
  assign mem_86_MPORT_1_addr = mem_86_MPORT_1_addr_pipe_0;
  assign mem_86_MPORT_1_data = mem_86[mem_86_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_86_MPORT_data = io_adcValues_86;
  assign mem_86_MPORT_addr = counter;
  assign mem_86_MPORT_mask = 1'h1;
  assign mem_86_MPORT_en = 1'h1;
  assign mem_87_MPORT_1_en = mem_87_MPORT_1_en_pipe_0;
  assign mem_87_MPORT_1_addr = mem_87_MPORT_1_addr_pipe_0;
  assign mem_87_MPORT_1_data = mem_87[mem_87_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_87_MPORT_data = io_adcValues_87;
  assign mem_87_MPORT_addr = counter;
  assign mem_87_MPORT_mask = 1'h1;
  assign mem_87_MPORT_en = 1'h1;
  assign mem_88_MPORT_1_en = mem_88_MPORT_1_en_pipe_0;
  assign mem_88_MPORT_1_addr = mem_88_MPORT_1_addr_pipe_0;
  assign mem_88_MPORT_1_data = mem_88[mem_88_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_88_MPORT_data = io_adcValues_88;
  assign mem_88_MPORT_addr = counter;
  assign mem_88_MPORT_mask = 1'h1;
  assign mem_88_MPORT_en = 1'h1;
  assign mem_89_MPORT_1_en = mem_89_MPORT_1_en_pipe_0;
  assign mem_89_MPORT_1_addr = mem_89_MPORT_1_addr_pipe_0;
  assign mem_89_MPORT_1_data = mem_89[mem_89_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_89_MPORT_data = io_adcValues_89;
  assign mem_89_MPORT_addr = counter;
  assign mem_89_MPORT_mask = 1'h1;
  assign mem_89_MPORT_en = 1'h1;
  assign mem_90_MPORT_1_en = mem_90_MPORT_1_en_pipe_0;
  assign mem_90_MPORT_1_addr = mem_90_MPORT_1_addr_pipe_0;
  assign mem_90_MPORT_1_data = mem_90[mem_90_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_90_MPORT_data = io_adcValues_90;
  assign mem_90_MPORT_addr = counter;
  assign mem_90_MPORT_mask = 1'h1;
  assign mem_90_MPORT_en = 1'h1;
  assign mem_91_MPORT_1_en = mem_91_MPORT_1_en_pipe_0;
  assign mem_91_MPORT_1_addr = mem_91_MPORT_1_addr_pipe_0;
  assign mem_91_MPORT_1_data = mem_91[mem_91_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_91_MPORT_data = io_adcValues_91;
  assign mem_91_MPORT_addr = counter;
  assign mem_91_MPORT_mask = 1'h1;
  assign mem_91_MPORT_en = 1'h1;
  assign mem_92_MPORT_1_en = mem_92_MPORT_1_en_pipe_0;
  assign mem_92_MPORT_1_addr = mem_92_MPORT_1_addr_pipe_0;
  assign mem_92_MPORT_1_data = mem_92[mem_92_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_92_MPORT_data = io_adcValues_92;
  assign mem_92_MPORT_addr = counter;
  assign mem_92_MPORT_mask = 1'h1;
  assign mem_92_MPORT_en = 1'h1;
  assign mem_93_MPORT_1_en = mem_93_MPORT_1_en_pipe_0;
  assign mem_93_MPORT_1_addr = mem_93_MPORT_1_addr_pipe_0;
  assign mem_93_MPORT_1_data = mem_93[mem_93_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_93_MPORT_data = io_adcValues_93;
  assign mem_93_MPORT_addr = counter;
  assign mem_93_MPORT_mask = 1'h1;
  assign mem_93_MPORT_en = 1'h1;
  assign mem_94_MPORT_1_en = mem_94_MPORT_1_en_pipe_0;
  assign mem_94_MPORT_1_addr = mem_94_MPORT_1_addr_pipe_0;
  assign mem_94_MPORT_1_data = mem_94[mem_94_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_94_MPORT_data = io_adcValues_94;
  assign mem_94_MPORT_addr = counter;
  assign mem_94_MPORT_mask = 1'h1;
  assign mem_94_MPORT_en = 1'h1;
  assign mem_95_MPORT_1_en = mem_95_MPORT_1_en_pipe_0;
  assign mem_95_MPORT_1_addr = mem_95_MPORT_1_addr_pipe_0;
  assign mem_95_MPORT_1_data = mem_95[mem_95_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_95_MPORT_data = io_adcValues_95;
  assign mem_95_MPORT_addr = counter;
  assign mem_95_MPORT_mask = 1'h1;
  assign mem_95_MPORT_en = 1'h1;
  assign mem_96_MPORT_1_en = mem_96_MPORT_1_en_pipe_0;
  assign mem_96_MPORT_1_addr = mem_96_MPORT_1_addr_pipe_0;
  assign mem_96_MPORT_1_data = mem_96[mem_96_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_96_MPORT_data = io_adcValues_96;
  assign mem_96_MPORT_addr = counter;
  assign mem_96_MPORT_mask = 1'h1;
  assign mem_96_MPORT_en = 1'h1;
  assign mem_97_MPORT_1_en = mem_97_MPORT_1_en_pipe_0;
  assign mem_97_MPORT_1_addr = mem_97_MPORT_1_addr_pipe_0;
  assign mem_97_MPORT_1_data = mem_97[mem_97_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_97_MPORT_data = io_adcValues_97;
  assign mem_97_MPORT_addr = counter;
  assign mem_97_MPORT_mask = 1'h1;
  assign mem_97_MPORT_en = 1'h1;
  assign mem_98_MPORT_1_en = mem_98_MPORT_1_en_pipe_0;
  assign mem_98_MPORT_1_addr = mem_98_MPORT_1_addr_pipe_0;
  assign mem_98_MPORT_1_data = mem_98[mem_98_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_98_MPORT_data = io_adcValues_98;
  assign mem_98_MPORT_addr = counter;
  assign mem_98_MPORT_mask = 1'h1;
  assign mem_98_MPORT_en = 1'h1;
  assign mem_99_MPORT_1_en = mem_99_MPORT_1_en_pipe_0;
  assign mem_99_MPORT_1_addr = mem_99_MPORT_1_addr_pipe_0;
  assign mem_99_MPORT_1_data = mem_99[mem_99_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_99_MPORT_data = io_adcValues_99;
  assign mem_99_MPORT_addr = counter;
  assign mem_99_MPORT_mask = 1'h1;
  assign mem_99_MPORT_en = 1'h1;
  assign mem_100_MPORT_1_en = mem_100_MPORT_1_en_pipe_0;
  assign mem_100_MPORT_1_addr = mem_100_MPORT_1_addr_pipe_0;
  assign mem_100_MPORT_1_data = mem_100[mem_100_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_100_MPORT_data = io_adcValues_100;
  assign mem_100_MPORT_addr = counter;
  assign mem_100_MPORT_mask = 1'h1;
  assign mem_100_MPORT_en = 1'h1;
  assign mem_101_MPORT_1_en = mem_101_MPORT_1_en_pipe_0;
  assign mem_101_MPORT_1_addr = mem_101_MPORT_1_addr_pipe_0;
  assign mem_101_MPORT_1_data = mem_101[mem_101_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_101_MPORT_data = io_adcValues_101;
  assign mem_101_MPORT_addr = counter;
  assign mem_101_MPORT_mask = 1'h1;
  assign mem_101_MPORT_en = 1'h1;
  assign mem_102_MPORT_1_en = mem_102_MPORT_1_en_pipe_0;
  assign mem_102_MPORT_1_addr = mem_102_MPORT_1_addr_pipe_0;
  assign mem_102_MPORT_1_data = mem_102[mem_102_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_102_MPORT_data = io_adcValues_102;
  assign mem_102_MPORT_addr = counter;
  assign mem_102_MPORT_mask = 1'h1;
  assign mem_102_MPORT_en = 1'h1;
  assign mem_103_MPORT_1_en = mem_103_MPORT_1_en_pipe_0;
  assign mem_103_MPORT_1_addr = mem_103_MPORT_1_addr_pipe_0;
  assign mem_103_MPORT_1_data = mem_103[mem_103_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_103_MPORT_data = io_adcValues_103;
  assign mem_103_MPORT_addr = counter;
  assign mem_103_MPORT_mask = 1'h1;
  assign mem_103_MPORT_en = 1'h1;
  assign mem_104_MPORT_1_en = mem_104_MPORT_1_en_pipe_0;
  assign mem_104_MPORT_1_addr = mem_104_MPORT_1_addr_pipe_0;
  assign mem_104_MPORT_1_data = mem_104[mem_104_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_104_MPORT_data = io_adcValues_104;
  assign mem_104_MPORT_addr = counter;
  assign mem_104_MPORT_mask = 1'h1;
  assign mem_104_MPORT_en = 1'h1;
  assign mem_105_MPORT_1_en = mem_105_MPORT_1_en_pipe_0;
  assign mem_105_MPORT_1_addr = mem_105_MPORT_1_addr_pipe_0;
  assign mem_105_MPORT_1_data = mem_105[mem_105_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_105_MPORT_data = io_adcValues_105;
  assign mem_105_MPORT_addr = counter;
  assign mem_105_MPORT_mask = 1'h1;
  assign mem_105_MPORT_en = 1'h1;
  assign mem_106_MPORT_1_en = mem_106_MPORT_1_en_pipe_0;
  assign mem_106_MPORT_1_addr = mem_106_MPORT_1_addr_pipe_0;
  assign mem_106_MPORT_1_data = mem_106[mem_106_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_106_MPORT_data = io_adcValues_106;
  assign mem_106_MPORT_addr = counter;
  assign mem_106_MPORT_mask = 1'h1;
  assign mem_106_MPORT_en = 1'h1;
  assign mem_107_MPORT_1_en = mem_107_MPORT_1_en_pipe_0;
  assign mem_107_MPORT_1_addr = mem_107_MPORT_1_addr_pipe_0;
  assign mem_107_MPORT_1_data = mem_107[mem_107_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_107_MPORT_data = io_adcValues_107;
  assign mem_107_MPORT_addr = counter;
  assign mem_107_MPORT_mask = 1'h1;
  assign mem_107_MPORT_en = 1'h1;
  assign mem_108_MPORT_1_en = mem_108_MPORT_1_en_pipe_0;
  assign mem_108_MPORT_1_addr = mem_108_MPORT_1_addr_pipe_0;
  assign mem_108_MPORT_1_data = mem_108[mem_108_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_108_MPORT_data = io_adcValues_108;
  assign mem_108_MPORT_addr = counter;
  assign mem_108_MPORT_mask = 1'h1;
  assign mem_108_MPORT_en = 1'h1;
  assign mem_109_MPORT_1_en = mem_109_MPORT_1_en_pipe_0;
  assign mem_109_MPORT_1_addr = mem_109_MPORT_1_addr_pipe_0;
  assign mem_109_MPORT_1_data = mem_109[mem_109_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_109_MPORT_data = io_adcValues_109;
  assign mem_109_MPORT_addr = counter;
  assign mem_109_MPORT_mask = 1'h1;
  assign mem_109_MPORT_en = 1'h1;
  assign mem_110_MPORT_1_en = mem_110_MPORT_1_en_pipe_0;
  assign mem_110_MPORT_1_addr = mem_110_MPORT_1_addr_pipe_0;
  assign mem_110_MPORT_1_data = mem_110[mem_110_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_110_MPORT_data = io_adcValues_110;
  assign mem_110_MPORT_addr = counter;
  assign mem_110_MPORT_mask = 1'h1;
  assign mem_110_MPORT_en = 1'h1;
  assign mem_111_MPORT_1_en = mem_111_MPORT_1_en_pipe_0;
  assign mem_111_MPORT_1_addr = mem_111_MPORT_1_addr_pipe_0;
  assign mem_111_MPORT_1_data = mem_111[mem_111_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_111_MPORT_data = io_adcValues_111;
  assign mem_111_MPORT_addr = counter;
  assign mem_111_MPORT_mask = 1'h1;
  assign mem_111_MPORT_en = 1'h1;
  assign mem_112_MPORT_1_en = mem_112_MPORT_1_en_pipe_0;
  assign mem_112_MPORT_1_addr = mem_112_MPORT_1_addr_pipe_0;
  assign mem_112_MPORT_1_data = mem_112[mem_112_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_112_MPORT_data = io_adcValues_112;
  assign mem_112_MPORT_addr = counter;
  assign mem_112_MPORT_mask = 1'h1;
  assign mem_112_MPORT_en = 1'h1;
  assign mem_113_MPORT_1_en = mem_113_MPORT_1_en_pipe_0;
  assign mem_113_MPORT_1_addr = mem_113_MPORT_1_addr_pipe_0;
  assign mem_113_MPORT_1_data = mem_113[mem_113_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_113_MPORT_data = io_adcValues_113;
  assign mem_113_MPORT_addr = counter;
  assign mem_113_MPORT_mask = 1'h1;
  assign mem_113_MPORT_en = 1'h1;
  assign mem_114_MPORT_1_en = mem_114_MPORT_1_en_pipe_0;
  assign mem_114_MPORT_1_addr = mem_114_MPORT_1_addr_pipe_0;
  assign mem_114_MPORT_1_data = mem_114[mem_114_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_114_MPORT_data = io_adcValues_114;
  assign mem_114_MPORT_addr = counter;
  assign mem_114_MPORT_mask = 1'h1;
  assign mem_114_MPORT_en = 1'h1;
  assign mem_115_MPORT_1_en = mem_115_MPORT_1_en_pipe_0;
  assign mem_115_MPORT_1_addr = mem_115_MPORT_1_addr_pipe_0;
  assign mem_115_MPORT_1_data = mem_115[mem_115_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_115_MPORT_data = io_adcValues_115;
  assign mem_115_MPORT_addr = counter;
  assign mem_115_MPORT_mask = 1'h1;
  assign mem_115_MPORT_en = 1'h1;
  assign mem_116_MPORT_1_en = mem_116_MPORT_1_en_pipe_0;
  assign mem_116_MPORT_1_addr = mem_116_MPORT_1_addr_pipe_0;
  assign mem_116_MPORT_1_data = mem_116[mem_116_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_116_MPORT_data = io_adcValues_116;
  assign mem_116_MPORT_addr = counter;
  assign mem_116_MPORT_mask = 1'h1;
  assign mem_116_MPORT_en = 1'h1;
  assign mem_117_MPORT_1_en = mem_117_MPORT_1_en_pipe_0;
  assign mem_117_MPORT_1_addr = mem_117_MPORT_1_addr_pipe_0;
  assign mem_117_MPORT_1_data = mem_117[mem_117_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_117_MPORT_data = io_adcValues_117;
  assign mem_117_MPORT_addr = counter;
  assign mem_117_MPORT_mask = 1'h1;
  assign mem_117_MPORT_en = 1'h1;
  assign mem_118_MPORT_1_en = mem_118_MPORT_1_en_pipe_0;
  assign mem_118_MPORT_1_addr = mem_118_MPORT_1_addr_pipe_0;
  assign mem_118_MPORT_1_data = mem_118[mem_118_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_118_MPORT_data = io_adcValues_118;
  assign mem_118_MPORT_addr = counter;
  assign mem_118_MPORT_mask = 1'h1;
  assign mem_118_MPORT_en = 1'h1;
  assign mem_119_MPORT_1_en = mem_119_MPORT_1_en_pipe_0;
  assign mem_119_MPORT_1_addr = mem_119_MPORT_1_addr_pipe_0;
  assign mem_119_MPORT_1_data = mem_119[mem_119_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_119_MPORT_data = io_adcValues_119;
  assign mem_119_MPORT_addr = counter;
  assign mem_119_MPORT_mask = 1'h1;
  assign mem_119_MPORT_en = 1'h1;
  assign mem_120_MPORT_1_en = mem_120_MPORT_1_en_pipe_0;
  assign mem_120_MPORT_1_addr = mem_120_MPORT_1_addr_pipe_0;
  assign mem_120_MPORT_1_data = mem_120[mem_120_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_120_MPORT_data = io_adcValues_120;
  assign mem_120_MPORT_addr = counter;
  assign mem_120_MPORT_mask = 1'h1;
  assign mem_120_MPORT_en = 1'h1;
  assign mem_121_MPORT_1_en = mem_121_MPORT_1_en_pipe_0;
  assign mem_121_MPORT_1_addr = mem_121_MPORT_1_addr_pipe_0;
  assign mem_121_MPORT_1_data = mem_121[mem_121_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_121_MPORT_data = io_adcValues_121;
  assign mem_121_MPORT_addr = counter;
  assign mem_121_MPORT_mask = 1'h1;
  assign mem_121_MPORT_en = 1'h1;
  assign mem_122_MPORT_1_en = mem_122_MPORT_1_en_pipe_0;
  assign mem_122_MPORT_1_addr = mem_122_MPORT_1_addr_pipe_0;
  assign mem_122_MPORT_1_data = mem_122[mem_122_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_122_MPORT_data = io_adcValues_122;
  assign mem_122_MPORT_addr = counter;
  assign mem_122_MPORT_mask = 1'h1;
  assign mem_122_MPORT_en = 1'h1;
  assign mem_123_MPORT_1_en = mem_123_MPORT_1_en_pipe_0;
  assign mem_123_MPORT_1_addr = mem_123_MPORT_1_addr_pipe_0;
  assign mem_123_MPORT_1_data = mem_123[mem_123_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_123_MPORT_data = io_adcValues_123;
  assign mem_123_MPORT_addr = counter;
  assign mem_123_MPORT_mask = 1'h1;
  assign mem_123_MPORT_en = 1'h1;
  assign mem_124_MPORT_1_en = mem_124_MPORT_1_en_pipe_0;
  assign mem_124_MPORT_1_addr = mem_124_MPORT_1_addr_pipe_0;
  assign mem_124_MPORT_1_data = mem_124[mem_124_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_124_MPORT_data = io_adcValues_124;
  assign mem_124_MPORT_addr = counter;
  assign mem_124_MPORT_mask = 1'h1;
  assign mem_124_MPORT_en = 1'h1;
  assign mem_125_MPORT_1_en = mem_125_MPORT_1_en_pipe_0;
  assign mem_125_MPORT_1_addr = mem_125_MPORT_1_addr_pipe_0;
  assign mem_125_MPORT_1_data = mem_125[mem_125_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_125_MPORT_data = io_adcValues_125;
  assign mem_125_MPORT_addr = counter;
  assign mem_125_MPORT_mask = 1'h1;
  assign mem_125_MPORT_en = 1'h1;
  assign mem_126_MPORT_1_en = mem_126_MPORT_1_en_pipe_0;
  assign mem_126_MPORT_1_addr = mem_126_MPORT_1_addr_pipe_0;
  assign mem_126_MPORT_1_data = mem_126[mem_126_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_126_MPORT_data = io_adcValues_126;
  assign mem_126_MPORT_addr = counter;
  assign mem_126_MPORT_mask = 1'h1;
  assign mem_126_MPORT_en = 1'h1;
  assign mem_127_MPORT_1_en = mem_127_MPORT_1_en_pipe_0;
  assign mem_127_MPORT_1_addr = mem_127_MPORT_1_addr_pipe_0;
  assign mem_127_MPORT_1_data = mem_127[mem_127_MPORT_1_addr]; // @[BufferMemorySystem.scala 16:24]
  assign mem_127_MPORT_data = io_adcValues_127;
  assign mem_127_MPORT_addr = counter;
  assign mem_127_MPORT_mask = 1'h1;
  assign mem_127_MPORT_en = 1'h1;
  assign io_dataOut_0 = mem_0_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_1 = mem_1_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_2 = mem_2_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_3 = mem_3_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_4 = mem_4_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_5 = mem_5_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_6 = mem_6_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_7 = mem_7_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_8 = mem_8_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_9 = mem_9_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_10 = mem_10_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_11 = mem_11_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_12 = mem_12_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_13 = mem_13_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_14 = mem_14_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_15 = mem_15_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_16 = mem_16_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_17 = mem_17_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_18 = mem_18_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_19 = mem_19_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_20 = mem_20_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_21 = mem_21_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_22 = mem_22_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_23 = mem_23_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_24 = mem_24_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_25 = mem_25_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_26 = mem_26_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_27 = mem_27_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_28 = mem_28_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_29 = mem_29_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_30 = mem_30_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_31 = mem_31_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_32 = mem_32_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_33 = mem_33_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_34 = mem_34_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_35 = mem_35_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_36 = mem_36_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_37 = mem_37_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_38 = mem_38_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_39 = mem_39_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_40 = mem_40_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_41 = mem_41_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_42 = mem_42_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_43 = mem_43_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_44 = mem_44_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_45 = mem_45_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_46 = mem_46_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_47 = mem_47_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_48 = mem_48_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_49 = mem_49_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_50 = mem_50_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_51 = mem_51_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_52 = mem_52_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_53 = mem_53_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_54 = mem_54_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_55 = mem_55_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_56 = mem_56_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_57 = mem_57_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_58 = mem_58_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_59 = mem_59_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_60 = mem_60_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_61 = mem_61_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_62 = mem_62_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_63 = mem_63_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_64 = mem_64_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_65 = mem_65_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_66 = mem_66_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_67 = mem_67_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_68 = mem_68_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_69 = mem_69_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_70 = mem_70_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_71 = mem_71_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_72 = mem_72_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_73 = mem_73_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_74 = mem_74_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_75 = mem_75_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_76 = mem_76_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_77 = mem_77_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_78 = mem_78_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_79 = mem_79_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_80 = mem_80_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_81 = mem_81_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_82 = mem_82_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_83 = mem_83_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_84 = mem_84_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_85 = mem_85_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_86 = mem_86_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_87 = mem_87_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_88 = mem_88_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_89 = mem_89_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_90 = mem_90_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_91 = mem_91_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_92 = mem_92_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_93 = mem_93_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_94 = mem_94_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_95 = mem_95_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_96 = mem_96_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_97 = mem_97_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_98 = mem_98_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_99 = mem_99_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_100 = mem_100_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_101 = mem_101_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_102 = mem_102_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_103 = mem_103_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_104 = mem_104_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_105 = mem_105_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_106 = mem_106_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_107 = mem_107_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_108 = mem_108_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_109 = mem_109_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_110 = mem_110_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_111 = mem_111_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_112 = mem_112_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_113 = mem_113_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_114 = mem_114_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_115 = mem_115_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_116 = mem_116_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_117 = mem_117_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_118 = mem_118_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_119 = mem_119_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_120 = mem_120_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_121 = mem_121_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_122 = mem_122_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_123 = mem_123_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_124 = mem_124_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_125 = mem_125_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_126 = mem_126_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  assign io_dataOut_127 = mem_127_MPORT_1_data; // @[BufferMemorySystem.scala 24:14]
  always @(posedge clock) begin
    if (mem_0_MPORT_en & mem_0_MPORT_mask) begin
      mem_0[mem_0_MPORT_addr] <= mem_0_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_0_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_0_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_1_MPORT_en & mem_1_MPORT_mask) begin
      mem_1[mem_1_MPORT_addr] <= mem_1_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_1_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_1_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_2_MPORT_en & mem_2_MPORT_mask) begin
      mem_2[mem_2_MPORT_addr] <= mem_2_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_2_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_2_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_3_MPORT_en & mem_3_MPORT_mask) begin
      mem_3[mem_3_MPORT_addr] <= mem_3_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_3_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_3_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_4_MPORT_en & mem_4_MPORT_mask) begin
      mem_4[mem_4_MPORT_addr] <= mem_4_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_4_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_4_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_5_MPORT_en & mem_5_MPORT_mask) begin
      mem_5[mem_5_MPORT_addr] <= mem_5_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_5_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_5_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_6_MPORT_en & mem_6_MPORT_mask) begin
      mem_6[mem_6_MPORT_addr] <= mem_6_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_6_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_6_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_7_MPORT_en & mem_7_MPORT_mask) begin
      mem_7[mem_7_MPORT_addr] <= mem_7_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_7_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_7_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_8_MPORT_en & mem_8_MPORT_mask) begin
      mem_8[mem_8_MPORT_addr] <= mem_8_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_8_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_8_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_9_MPORT_en & mem_9_MPORT_mask) begin
      mem_9[mem_9_MPORT_addr] <= mem_9_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_9_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_9_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_10_MPORT_en & mem_10_MPORT_mask) begin
      mem_10[mem_10_MPORT_addr] <= mem_10_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_10_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_10_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_11_MPORT_en & mem_11_MPORT_mask) begin
      mem_11[mem_11_MPORT_addr] <= mem_11_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_11_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_11_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_12_MPORT_en & mem_12_MPORT_mask) begin
      mem_12[mem_12_MPORT_addr] <= mem_12_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_12_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_12_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_13_MPORT_en & mem_13_MPORT_mask) begin
      mem_13[mem_13_MPORT_addr] <= mem_13_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_13_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_13_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_14_MPORT_en & mem_14_MPORT_mask) begin
      mem_14[mem_14_MPORT_addr] <= mem_14_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_14_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_14_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_15_MPORT_en & mem_15_MPORT_mask) begin
      mem_15[mem_15_MPORT_addr] <= mem_15_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_15_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_15_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_16_MPORT_en & mem_16_MPORT_mask) begin
      mem_16[mem_16_MPORT_addr] <= mem_16_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_16_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_16_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_17_MPORT_en & mem_17_MPORT_mask) begin
      mem_17[mem_17_MPORT_addr] <= mem_17_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_17_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_17_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_18_MPORT_en & mem_18_MPORT_mask) begin
      mem_18[mem_18_MPORT_addr] <= mem_18_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_18_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_18_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_19_MPORT_en & mem_19_MPORT_mask) begin
      mem_19[mem_19_MPORT_addr] <= mem_19_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_19_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_19_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_20_MPORT_en & mem_20_MPORT_mask) begin
      mem_20[mem_20_MPORT_addr] <= mem_20_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_20_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_20_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_21_MPORT_en & mem_21_MPORT_mask) begin
      mem_21[mem_21_MPORT_addr] <= mem_21_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_21_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_21_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_22_MPORT_en & mem_22_MPORT_mask) begin
      mem_22[mem_22_MPORT_addr] <= mem_22_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_22_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_22_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_23_MPORT_en & mem_23_MPORT_mask) begin
      mem_23[mem_23_MPORT_addr] <= mem_23_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_23_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_23_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_24_MPORT_en & mem_24_MPORT_mask) begin
      mem_24[mem_24_MPORT_addr] <= mem_24_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_24_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_24_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_25_MPORT_en & mem_25_MPORT_mask) begin
      mem_25[mem_25_MPORT_addr] <= mem_25_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_25_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_25_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_26_MPORT_en & mem_26_MPORT_mask) begin
      mem_26[mem_26_MPORT_addr] <= mem_26_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_26_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_26_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_27_MPORT_en & mem_27_MPORT_mask) begin
      mem_27[mem_27_MPORT_addr] <= mem_27_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_27_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_27_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_28_MPORT_en & mem_28_MPORT_mask) begin
      mem_28[mem_28_MPORT_addr] <= mem_28_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_28_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_28_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_29_MPORT_en & mem_29_MPORT_mask) begin
      mem_29[mem_29_MPORT_addr] <= mem_29_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_29_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_29_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_30_MPORT_en & mem_30_MPORT_mask) begin
      mem_30[mem_30_MPORT_addr] <= mem_30_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_30_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_30_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_31_MPORT_en & mem_31_MPORT_mask) begin
      mem_31[mem_31_MPORT_addr] <= mem_31_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_31_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_31_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_32_MPORT_en & mem_32_MPORT_mask) begin
      mem_32[mem_32_MPORT_addr] <= mem_32_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_32_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_32_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_33_MPORT_en & mem_33_MPORT_mask) begin
      mem_33[mem_33_MPORT_addr] <= mem_33_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_33_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_33_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_34_MPORT_en & mem_34_MPORT_mask) begin
      mem_34[mem_34_MPORT_addr] <= mem_34_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_34_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_34_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_35_MPORT_en & mem_35_MPORT_mask) begin
      mem_35[mem_35_MPORT_addr] <= mem_35_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_35_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_35_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_36_MPORT_en & mem_36_MPORT_mask) begin
      mem_36[mem_36_MPORT_addr] <= mem_36_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_36_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_36_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_37_MPORT_en & mem_37_MPORT_mask) begin
      mem_37[mem_37_MPORT_addr] <= mem_37_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_37_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_37_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_38_MPORT_en & mem_38_MPORT_mask) begin
      mem_38[mem_38_MPORT_addr] <= mem_38_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_38_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_38_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_39_MPORT_en & mem_39_MPORT_mask) begin
      mem_39[mem_39_MPORT_addr] <= mem_39_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_39_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_39_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_40_MPORT_en & mem_40_MPORT_mask) begin
      mem_40[mem_40_MPORT_addr] <= mem_40_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_40_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_40_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_41_MPORT_en & mem_41_MPORT_mask) begin
      mem_41[mem_41_MPORT_addr] <= mem_41_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_41_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_41_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_42_MPORT_en & mem_42_MPORT_mask) begin
      mem_42[mem_42_MPORT_addr] <= mem_42_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_42_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_42_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_43_MPORT_en & mem_43_MPORT_mask) begin
      mem_43[mem_43_MPORT_addr] <= mem_43_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_43_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_43_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_44_MPORT_en & mem_44_MPORT_mask) begin
      mem_44[mem_44_MPORT_addr] <= mem_44_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_44_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_44_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_45_MPORT_en & mem_45_MPORT_mask) begin
      mem_45[mem_45_MPORT_addr] <= mem_45_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_45_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_45_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_46_MPORT_en & mem_46_MPORT_mask) begin
      mem_46[mem_46_MPORT_addr] <= mem_46_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_46_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_46_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_47_MPORT_en & mem_47_MPORT_mask) begin
      mem_47[mem_47_MPORT_addr] <= mem_47_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_47_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_47_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_48_MPORT_en & mem_48_MPORT_mask) begin
      mem_48[mem_48_MPORT_addr] <= mem_48_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_48_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_48_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_49_MPORT_en & mem_49_MPORT_mask) begin
      mem_49[mem_49_MPORT_addr] <= mem_49_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_49_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_49_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_50_MPORT_en & mem_50_MPORT_mask) begin
      mem_50[mem_50_MPORT_addr] <= mem_50_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_50_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_50_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_51_MPORT_en & mem_51_MPORT_mask) begin
      mem_51[mem_51_MPORT_addr] <= mem_51_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_51_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_51_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_52_MPORT_en & mem_52_MPORT_mask) begin
      mem_52[mem_52_MPORT_addr] <= mem_52_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_52_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_52_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_53_MPORT_en & mem_53_MPORT_mask) begin
      mem_53[mem_53_MPORT_addr] <= mem_53_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_53_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_53_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_54_MPORT_en & mem_54_MPORT_mask) begin
      mem_54[mem_54_MPORT_addr] <= mem_54_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_54_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_54_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_55_MPORT_en & mem_55_MPORT_mask) begin
      mem_55[mem_55_MPORT_addr] <= mem_55_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_55_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_55_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_56_MPORT_en & mem_56_MPORT_mask) begin
      mem_56[mem_56_MPORT_addr] <= mem_56_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_56_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_56_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_57_MPORT_en & mem_57_MPORT_mask) begin
      mem_57[mem_57_MPORT_addr] <= mem_57_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_57_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_57_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_58_MPORT_en & mem_58_MPORT_mask) begin
      mem_58[mem_58_MPORT_addr] <= mem_58_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_58_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_58_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_59_MPORT_en & mem_59_MPORT_mask) begin
      mem_59[mem_59_MPORT_addr] <= mem_59_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_59_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_59_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_60_MPORT_en & mem_60_MPORT_mask) begin
      mem_60[mem_60_MPORT_addr] <= mem_60_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_60_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_60_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_61_MPORT_en & mem_61_MPORT_mask) begin
      mem_61[mem_61_MPORT_addr] <= mem_61_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_61_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_61_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_62_MPORT_en & mem_62_MPORT_mask) begin
      mem_62[mem_62_MPORT_addr] <= mem_62_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_62_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_62_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_63_MPORT_en & mem_63_MPORT_mask) begin
      mem_63[mem_63_MPORT_addr] <= mem_63_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_63_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_63_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_64_MPORT_en & mem_64_MPORT_mask) begin
      mem_64[mem_64_MPORT_addr] <= mem_64_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_64_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_64_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_65_MPORT_en & mem_65_MPORT_mask) begin
      mem_65[mem_65_MPORT_addr] <= mem_65_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_65_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_65_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_66_MPORT_en & mem_66_MPORT_mask) begin
      mem_66[mem_66_MPORT_addr] <= mem_66_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_66_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_66_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_67_MPORT_en & mem_67_MPORT_mask) begin
      mem_67[mem_67_MPORT_addr] <= mem_67_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_67_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_67_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_68_MPORT_en & mem_68_MPORT_mask) begin
      mem_68[mem_68_MPORT_addr] <= mem_68_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_68_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_68_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_69_MPORT_en & mem_69_MPORT_mask) begin
      mem_69[mem_69_MPORT_addr] <= mem_69_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_69_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_69_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_70_MPORT_en & mem_70_MPORT_mask) begin
      mem_70[mem_70_MPORT_addr] <= mem_70_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_70_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_70_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_71_MPORT_en & mem_71_MPORT_mask) begin
      mem_71[mem_71_MPORT_addr] <= mem_71_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_71_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_71_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_72_MPORT_en & mem_72_MPORT_mask) begin
      mem_72[mem_72_MPORT_addr] <= mem_72_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_72_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_72_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_73_MPORT_en & mem_73_MPORT_mask) begin
      mem_73[mem_73_MPORT_addr] <= mem_73_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_73_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_73_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_74_MPORT_en & mem_74_MPORT_mask) begin
      mem_74[mem_74_MPORT_addr] <= mem_74_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_74_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_74_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_75_MPORT_en & mem_75_MPORT_mask) begin
      mem_75[mem_75_MPORT_addr] <= mem_75_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_75_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_75_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_76_MPORT_en & mem_76_MPORT_mask) begin
      mem_76[mem_76_MPORT_addr] <= mem_76_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_76_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_76_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_77_MPORT_en & mem_77_MPORT_mask) begin
      mem_77[mem_77_MPORT_addr] <= mem_77_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_77_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_77_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_78_MPORT_en & mem_78_MPORT_mask) begin
      mem_78[mem_78_MPORT_addr] <= mem_78_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_78_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_78_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_79_MPORT_en & mem_79_MPORT_mask) begin
      mem_79[mem_79_MPORT_addr] <= mem_79_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_79_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_79_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_80_MPORT_en & mem_80_MPORT_mask) begin
      mem_80[mem_80_MPORT_addr] <= mem_80_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_80_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_80_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_81_MPORT_en & mem_81_MPORT_mask) begin
      mem_81[mem_81_MPORT_addr] <= mem_81_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_81_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_81_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_82_MPORT_en & mem_82_MPORT_mask) begin
      mem_82[mem_82_MPORT_addr] <= mem_82_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_82_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_82_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_83_MPORT_en & mem_83_MPORT_mask) begin
      mem_83[mem_83_MPORT_addr] <= mem_83_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_83_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_83_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_84_MPORT_en & mem_84_MPORT_mask) begin
      mem_84[mem_84_MPORT_addr] <= mem_84_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_84_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_84_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_85_MPORT_en & mem_85_MPORT_mask) begin
      mem_85[mem_85_MPORT_addr] <= mem_85_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_85_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_85_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_86_MPORT_en & mem_86_MPORT_mask) begin
      mem_86[mem_86_MPORT_addr] <= mem_86_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_86_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_86_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_87_MPORT_en & mem_87_MPORT_mask) begin
      mem_87[mem_87_MPORT_addr] <= mem_87_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_87_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_87_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_88_MPORT_en & mem_88_MPORT_mask) begin
      mem_88[mem_88_MPORT_addr] <= mem_88_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_88_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_88_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_89_MPORT_en & mem_89_MPORT_mask) begin
      mem_89[mem_89_MPORT_addr] <= mem_89_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_89_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_89_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_90_MPORT_en & mem_90_MPORT_mask) begin
      mem_90[mem_90_MPORT_addr] <= mem_90_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_90_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_90_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_91_MPORT_en & mem_91_MPORT_mask) begin
      mem_91[mem_91_MPORT_addr] <= mem_91_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_91_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_91_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_92_MPORT_en & mem_92_MPORT_mask) begin
      mem_92[mem_92_MPORT_addr] <= mem_92_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_92_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_92_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_93_MPORT_en & mem_93_MPORT_mask) begin
      mem_93[mem_93_MPORT_addr] <= mem_93_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_93_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_93_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_94_MPORT_en & mem_94_MPORT_mask) begin
      mem_94[mem_94_MPORT_addr] <= mem_94_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_94_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_94_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_95_MPORT_en & mem_95_MPORT_mask) begin
      mem_95[mem_95_MPORT_addr] <= mem_95_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_95_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_95_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_96_MPORT_en & mem_96_MPORT_mask) begin
      mem_96[mem_96_MPORT_addr] <= mem_96_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_96_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_96_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_97_MPORT_en & mem_97_MPORT_mask) begin
      mem_97[mem_97_MPORT_addr] <= mem_97_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_97_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_97_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_98_MPORT_en & mem_98_MPORT_mask) begin
      mem_98[mem_98_MPORT_addr] <= mem_98_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_98_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_98_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_99_MPORT_en & mem_99_MPORT_mask) begin
      mem_99[mem_99_MPORT_addr] <= mem_99_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_99_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_99_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_100_MPORT_en & mem_100_MPORT_mask) begin
      mem_100[mem_100_MPORT_addr] <= mem_100_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_100_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_100_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_101_MPORT_en & mem_101_MPORT_mask) begin
      mem_101[mem_101_MPORT_addr] <= mem_101_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_101_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_101_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_102_MPORT_en & mem_102_MPORT_mask) begin
      mem_102[mem_102_MPORT_addr] <= mem_102_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_102_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_102_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_103_MPORT_en & mem_103_MPORT_mask) begin
      mem_103[mem_103_MPORT_addr] <= mem_103_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_103_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_103_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_104_MPORT_en & mem_104_MPORT_mask) begin
      mem_104[mem_104_MPORT_addr] <= mem_104_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_104_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_104_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_105_MPORT_en & mem_105_MPORT_mask) begin
      mem_105[mem_105_MPORT_addr] <= mem_105_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_105_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_105_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_106_MPORT_en & mem_106_MPORT_mask) begin
      mem_106[mem_106_MPORT_addr] <= mem_106_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_106_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_106_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_107_MPORT_en & mem_107_MPORT_mask) begin
      mem_107[mem_107_MPORT_addr] <= mem_107_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_107_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_107_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_108_MPORT_en & mem_108_MPORT_mask) begin
      mem_108[mem_108_MPORT_addr] <= mem_108_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_108_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_108_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_109_MPORT_en & mem_109_MPORT_mask) begin
      mem_109[mem_109_MPORT_addr] <= mem_109_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_109_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_109_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_110_MPORT_en & mem_110_MPORT_mask) begin
      mem_110[mem_110_MPORT_addr] <= mem_110_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_110_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_110_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_111_MPORT_en & mem_111_MPORT_mask) begin
      mem_111[mem_111_MPORT_addr] <= mem_111_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_111_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_111_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_112_MPORT_en & mem_112_MPORT_mask) begin
      mem_112[mem_112_MPORT_addr] <= mem_112_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_112_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_112_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_113_MPORT_en & mem_113_MPORT_mask) begin
      mem_113[mem_113_MPORT_addr] <= mem_113_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_113_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_113_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_114_MPORT_en & mem_114_MPORT_mask) begin
      mem_114[mem_114_MPORT_addr] <= mem_114_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_114_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_114_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_115_MPORT_en & mem_115_MPORT_mask) begin
      mem_115[mem_115_MPORT_addr] <= mem_115_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_115_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_115_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_116_MPORT_en & mem_116_MPORT_mask) begin
      mem_116[mem_116_MPORT_addr] <= mem_116_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_116_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_116_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_117_MPORT_en & mem_117_MPORT_mask) begin
      mem_117[mem_117_MPORT_addr] <= mem_117_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_117_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_117_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_118_MPORT_en & mem_118_MPORT_mask) begin
      mem_118[mem_118_MPORT_addr] <= mem_118_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_118_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_118_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_119_MPORT_en & mem_119_MPORT_mask) begin
      mem_119[mem_119_MPORT_addr] <= mem_119_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_119_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_119_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_120_MPORT_en & mem_120_MPORT_mask) begin
      mem_120[mem_120_MPORT_addr] <= mem_120_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_120_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_120_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_121_MPORT_en & mem_121_MPORT_mask) begin
      mem_121[mem_121_MPORT_addr] <= mem_121_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_121_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_121_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_122_MPORT_en & mem_122_MPORT_mask) begin
      mem_122[mem_122_MPORT_addr] <= mem_122_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_122_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_122_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_123_MPORT_en & mem_123_MPORT_mask) begin
      mem_123[mem_123_MPORT_addr] <= mem_123_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_123_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_123_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_124_MPORT_en & mem_124_MPORT_mask) begin
      mem_124[mem_124_MPORT_addr] <= mem_124_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_124_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_124_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_125_MPORT_en & mem_125_MPORT_mask) begin
      mem_125[mem_125_MPORT_addr] <= mem_125_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_125_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_125_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_126_MPORT_en & mem_126_MPORT_mask) begin
      mem_126[mem_126_MPORT_addr] <= mem_126_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_126_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_126_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (mem_127_MPORT_en & mem_127_MPORT_mask) begin
      mem_127[mem_127_MPORT_addr] <= mem_127_MPORT_data; // @[BufferMemorySystem.scala 16:24]
    end
    mem_127_MPORT_1_en_pipe_0 <= io_enable;
    if (io_enable) begin
      mem_127_MPORT_1_addr_pipe_0 <= io_addr;
    end
    if (reset) begin // @[BufferMemorySystem.scala 14:24]
      counter <= 4'h0; // @[BufferMemorySystem.scala 14:24]
    end else if (io_enable) begin // @[BufferMemorySystem.scala 18:39]
      counter <= _counter_T_1; // @[BufferMemorySystem.scala 19:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_0[initvar] = _RAND_0[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_1[initvar] = _RAND_3[7:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_2[initvar] = _RAND_6[7:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_3[initvar] = _RAND_9[7:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_4[initvar] = _RAND_12[7:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_5[initvar] = _RAND_15[7:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_6[initvar] = _RAND_18[7:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_7[initvar] = _RAND_21[7:0];
  _RAND_24 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_8[initvar] = _RAND_24[7:0];
  _RAND_27 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_9[initvar] = _RAND_27[7:0];
  _RAND_30 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_10[initvar] = _RAND_30[7:0];
  _RAND_33 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_11[initvar] = _RAND_33[7:0];
  _RAND_36 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_12[initvar] = _RAND_36[7:0];
  _RAND_39 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_13[initvar] = _RAND_39[7:0];
  _RAND_42 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_14[initvar] = _RAND_42[7:0];
  _RAND_45 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_15[initvar] = _RAND_45[7:0];
  _RAND_48 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_16[initvar] = _RAND_48[7:0];
  _RAND_51 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_17[initvar] = _RAND_51[7:0];
  _RAND_54 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_18[initvar] = _RAND_54[7:0];
  _RAND_57 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_19[initvar] = _RAND_57[7:0];
  _RAND_60 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_20[initvar] = _RAND_60[7:0];
  _RAND_63 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_21[initvar] = _RAND_63[7:0];
  _RAND_66 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_22[initvar] = _RAND_66[7:0];
  _RAND_69 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_23[initvar] = _RAND_69[7:0];
  _RAND_72 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_24[initvar] = _RAND_72[7:0];
  _RAND_75 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_25[initvar] = _RAND_75[7:0];
  _RAND_78 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_26[initvar] = _RAND_78[7:0];
  _RAND_81 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_27[initvar] = _RAND_81[7:0];
  _RAND_84 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_28[initvar] = _RAND_84[7:0];
  _RAND_87 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_29[initvar] = _RAND_87[7:0];
  _RAND_90 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_30[initvar] = _RAND_90[7:0];
  _RAND_93 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_31[initvar] = _RAND_93[7:0];
  _RAND_96 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_32[initvar] = _RAND_96[7:0];
  _RAND_99 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_33[initvar] = _RAND_99[7:0];
  _RAND_102 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_34[initvar] = _RAND_102[7:0];
  _RAND_105 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_35[initvar] = _RAND_105[7:0];
  _RAND_108 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_36[initvar] = _RAND_108[7:0];
  _RAND_111 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_37[initvar] = _RAND_111[7:0];
  _RAND_114 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_38[initvar] = _RAND_114[7:0];
  _RAND_117 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_39[initvar] = _RAND_117[7:0];
  _RAND_120 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_40[initvar] = _RAND_120[7:0];
  _RAND_123 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_41[initvar] = _RAND_123[7:0];
  _RAND_126 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_42[initvar] = _RAND_126[7:0];
  _RAND_129 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_43[initvar] = _RAND_129[7:0];
  _RAND_132 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_44[initvar] = _RAND_132[7:0];
  _RAND_135 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_45[initvar] = _RAND_135[7:0];
  _RAND_138 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_46[initvar] = _RAND_138[7:0];
  _RAND_141 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_47[initvar] = _RAND_141[7:0];
  _RAND_144 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_48[initvar] = _RAND_144[7:0];
  _RAND_147 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_49[initvar] = _RAND_147[7:0];
  _RAND_150 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_50[initvar] = _RAND_150[7:0];
  _RAND_153 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_51[initvar] = _RAND_153[7:0];
  _RAND_156 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_52[initvar] = _RAND_156[7:0];
  _RAND_159 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_53[initvar] = _RAND_159[7:0];
  _RAND_162 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_54[initvar] = _RAND_162[7:0];
  _RAND_165 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_55[initvar] = _RAND_165[7:0];
  _RAND_168 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_56[initvar] = _RAND_168[7:0];
  _RAND_171 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_57[initvar] = _RAND_171[7:0];
  _RAND_174 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_58[initvar] = _RAND_174[7:0];
  _RAND_177 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_59[initvar] = _RAND_177[7:0];
  _RAND_180 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_60[initvar] = _RAND_180[7:0];
  _RAND_183 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_61[initvar] = _RAND_183[7:0];
  _RAND_186 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_62[initvar] = _RAND_186[7:0];
  _RAND_189 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_63[initvar] = _RAND_189[7:0];
  _RAND_192 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_64[initvar] = _RAND_192[7:0];
  _RAND_195 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_65[initvar] = _RAND_195[7:0];
  _RAND_198 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_66[initvar] = _RAND_198[7:0];
  _RAND_201 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_67[initvar] = _RAND_201[7:0];
  _RAND_204 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_68[initvar] = _RAND_204[7:0];
  _RAND_207 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_69[initvar] = _RAND_207[7:0];
  _RAND_210 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_70[initvar] = _RAND_210[7:0];
  _RAND_213 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_71[initvar] = _RAND_213[7:0];
  _RAND_216 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_72[initvar] = _RAND_216[7:0];
  _RAND_219 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_73[initvar] = _RAND_219[7:0];
  _RAND_222 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_74[initvar] = _RAND_222[7:0];
  _RAND_225 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_75[initvar] = _RAND_225[7:0];
  _RAND_228 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_76[initvar] = _RAND_228[7:0];
  _RAND_231 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_77[initvar] = _RAND_231[7:0];
  _RAND_234 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_78[initvar] = _RAND_234[7:0];
  _RAND_237 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_79[initvar] = _RAND_237[7:0];
  _RAND_240 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_80[initvar] = _RAND_240[7:0];
  _RAND_243 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_81[initvar] = _RAND_243[7:0];
  _RAND_246 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_82[initvar] = _RAND_246[7:0];
  _RAND_249 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_83[initvar] = _RAND_249[7:0];
  _RAND_252 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_84[initvar] = _RAND_252[7:0];
  _RAND_255 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_85[initvar] = _RAND_255[7:0];
  _RAND_258 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_86[initvar] = _RAND_258[7:0];
  _RAND_261 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_87[initvar] = _RAND_261[7:0];
  _RAND_264 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_88[initvar] = _RAND_264[7:0];
  _RAND_267 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_89[initvar] = _RAND_267[7:0];
  _RAND_270 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_90[initvar] = _RAND_270[7:0];
  _RAND_273 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_91[initvar] = _RAND_273[7:0];
  _RAND_276 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_92[initvar] = _RAND_276[7:0];
  _RAND_279 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_93[initvar] = _RAND_279[7:0];
  _RAND_282 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_94[initvar] = _RAND_282[7:0];
  _RAND_285 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_95[initvar] = _RAND_285[7:0];
  _RAND_288 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_96[initvar] = _RAND_288[7:0];
  _RAND_291 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_97[initvar] = _RAND_291[7:0];
  _RAND_294 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_98[initvar] = _RAND_294[7:0];
  _RAND_297 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_99[initvar] = _RAND_297[7:0];
  _RAND_300 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_100[initvar] = _RAND_300[7:0];
  _RAND_303 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_101[initvar] = _RAND_303[7:0];
  _RAND_306 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_102[initvar] = _RAND_306[7:0];
  _RAND_309 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_103[initvar] = _RAND_309[7:0];
  _RAND_312 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_104[initvar] = _RAND_312[7:0];
  _RAND_315 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_105[initvar] = _RAND_315[7:0];
  _RAND_318 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_106[initvar] = _RAND_318[7:0];
  _RAND_321 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_107[initvar] = _RAND_321[7:0];
  _RAND_324 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_108[initvar] = _RAND_324[7:0];
  _RAND_327 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_109[initvar] = _RAND_327[7:0];
  _RAND_330 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_110[initvar] = _RAND_330[7:0];
  _RAND_333 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_111[initvar] = _RAND_333[7:0];
  _RAND_336 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_112[initvar] = _RAND_336[7:0];
  _RAND_339 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_113[initvar] = _RAND_339[7:0];
  _RAND_342 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_114[initvar] = _RAND_342[7:0];
  _RAND_345 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_115[initvar] = _RAND_345[7:0];
  _RAND_348 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_116[initvar] = _RAND_348[7:0];
  _RAND_351 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_117[initvar] = _RAND_351[7:0];
  _RAND_354 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_118[initvar] = _RAND_354[7:0];
  _RAND_357 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_119[initvar] = _RAND_357[7:0];
  _RAND_360 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_120[initvar] = _RAND_360[7:0];
  _RAND_363 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_121[initvar] = _RAND_363[7:0];
  _RAND_366 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_122[initvar] = _RAND_366[7:0];
  _RAND_369 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_123[initvar] = _RAND_369[7:0];
  _RAND_372 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_124[initvar] = _RAND_372[7:0];
  _RAND_375 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_125[initvar] = _RAND_375[7:0];
  _RAND_378 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_126[initvar] = _RAND_378[7:0];
  _RAND_381 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mem_127[initvar] = _RAND_381[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_0_MPORT_1_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_0_MPORT_1_addr_pipe_0 = _RAND_2[3:0];
  _RAND_4 = {1{`RANDOM}};
  mem_1_MPORT_1_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  mem_1_MPORT_1_addr_pipe_0 = _RAND_5[3:0];
  _RAND_7 = {1{`RANDOM}};
  mem_2_MPORT_1_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  mem_2_MPORT_1_addr_pipe_0 = _RAND_8[3:0];
  _RAND_10 = {1{`RANDOM}};
  mem_3_MPORT_1_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  mem_3_MPORT_1_addr_pipe_0 = _RAND_11[3:0];
  _RAND_13 = {1{`RANDOM}};
  mem_4_MPORT_1_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  mem_4_MPORT_1_addr_pipe_0 = _RAND_14[3:0];
  _RAND_16 = {1{`RANDOM}};
  mem_5_MPORT_1_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  mem_5_MPORT_1_addr_pipe_0 = _RAND_17[3:0];
  _RAND_19 = {1{`RANDOM}};
  mem_6_MPORT_1_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  mem_6_MPORT_1_addr_pipe_0 = _RAND_20[3:0];
  _RAND_22 = {1{`RANDOM}};
  mem_7_MPORT_1_en_pipe_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  mem_7_MPORT_1_addr_pipe_0 = _RAND_23[3:0];
  _RAND_25 = {1{`RANDOM}};
  mem_8_MPORT_1_en_pipe_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  mem_8_MPORT_1_addr_pipe_0 = _RAND_26[3:0];
  _RAND_28 = {1{`RANDOM}};
  mem_9_MPORT_1_en_pipe_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  mem_9_MPORT_1_addr_pipe_0 = _RAND_29[3:0];
  _RAND_31 = {1{`RANDOM}};
  mem_10_MPORT_1_en_pipe_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  mem_10_MPORT_1_addr_pipe_0 = _RAND_32[3:0];
  _RAND_34 = {1{`RANDOM}};
  mem_11_MPORT_1_en_pipe_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  mem_11_MPORT_1_addr_pipe_0 = _RAND_35[3:0];
  _RAND_37 = {1{`RANDOM}};
  mem_12_MPORT_1_en_pipe_0 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  mem_12_MPORT_1_addr_pipe_0 = _RAND_38[3:0];
  _RAND_40 = {1{`RANDOM}};
  mem_13_MPORT_1_en_pipe_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  mem_13_MPORT_1_addr_pipe_0 = _RAND_41[3:0];
  _RAND_43 = {1{`RANDOM}};
  mem_14_MPORT_1_en_pipe_0 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  mem_14_MPORT_1_addr_pipe_0 = _RAND_44[3:0];
  _RAND_46 = {1{`RANDOM}};
  mem_15_MPORT_1_en_pipe_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  mem_15_MPORT_1_addr_pipe_0 = _RAND_47[3:0];
  _RAND_49 = {1{`RANDOM}};
  mem_16_MPORT_1_en_pipe_0 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  mem_16_MPORT_1_addr_pipe_0 = _RAND_50[3:0];
  _RAND_52 = {1{`RANDOM}};
  mem_17_MPORT_1_en_pipe_0 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  mem_17_MPORT_1_addr_pipe_0 = _RAND_53[3:0];
  _RAND_55 = {1{`RANDOM}};
  mem_18_MPORT_1_en_pipe_0 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  mem_18_MPORT_1_addr_pipe_0 = _RAND_56[3:0];
  _RAND_58 = {1{`RANDOM}};
  mem_19_MPORT_1_en_pipe_0 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  mem_19_MPORT_1_addr_pipe_0 = _RAND_59[3:0];
  _RAND_61 = {1{`RANDOM}};
  mem_20_MPORT_1_en_pipe_0 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  mem_20_MPORT_1_addr_pipe_0 = _RAND_62[3:0];
  _RAND_64 = {1{`RANDOM}};
  mem_21_MPORT_1_en_pipe_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  mem_21_MPORT_1_addr_pipe_0 = _RAND_65[3:0];
  _RAND_67 = {1{`RANDOM}};
  mem_22_MPORT_1_en_pipe_0 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  mem_22_MPORT_1_addr_pipe_0 = _RAND_68[3:0];
  _RAND_70 = {1{`RANDOM}};
  mem_23_MPORT_1_en_pipe_0 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  mem_23_MPORT_1_addr_pipe_0 = _RAND_71[3:0];
  _RAND_73 = {1{`RANDOM}};
  mem_24_MPORT_1_en_pipe_0 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  mem_24_MPORT_1_addr_pipe_0 = _RAND_74[3:0];
  _RAND_76 = {1{`RANDOM}};
  mem_25_MPORT_1_en_pipe_0 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  mem_25_MPORT_1_addr_pipe_0 = _RAND_77[3:0];
  _RAND_79 = {1{`RANDOM}};
  mem_26_MPORT_1_en_pipe_0 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  mem_26_MPORT_1_addr_pipe_0 = _RAND_80[3:0];
  _RAND_82 = {1{`RANDOM}};
  mem_27_MPORT_1_en_pipe_0 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  mem_27_MPORT_1_addr_pipe_0 = _RAND_83[3:0];
  _RAND_85 = {1{`RANDOM}};
  mem_28_MPORT_1_en_pipe_0 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  mem_28_MPORT_1_addr_pipe_0 = _RAND_86[3:0];
  _RAND_88 = {1{`RANDOM}};
  mem_29_MPORT_1_en_pipe_0 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  mem_29_MPORT_1_addr_pipe_0 = _RAND_89[3:0];
  _RAND_91 = {1{`RANDOM}};
  mem_30_MPORT_1_en_pipe_0 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  mem_30_MPORT_1_addr_pipe_0 = _RAND_92[3:0];
  _RAND_94 = {1{`RANDOM}};
  mem_31_MPORT_1_en_pipe_0 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  mem_31_MPORT_1_addr_pipe_0 = _RAND_95[3:0];
  _RAND_97 = {1{`RANDOM}};
  mem_32_MPORT_1_en_pipe_0 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  mem_32_MPORT_1_addr_pipe_0 = _RAND_98[3:0];
  _RAND_100 = {1{`RANDOM}};
  mem_33_MPORT_1_en_pipe_0 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  mem_33_MPORT_1_addr_pipe_0 = _RAND_101[3:0];
  _RAND_103 = {1{`RANDOM}};
  mem_34_MPORT_1_en_pipe_0 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  mem_34_MPORT_1_addr_pipe_0 = _RAND_104[3:0];
  _RAND_106 = {1{`RANDOM}};
  mem_35_MPORT_1_en_pipe_0 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  mem_35_MPORT_1_addr_pipe_0 = _RAND_107[3:0];
  _RAND_109 = {1{`RANDOM}};
  mem_36_MPORT_1_en_pipe_0 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  mem_36_MPORT_1_addr_pipe_0 = _RAND_110[3:0];
  _RAND_112 = {1{`RANDOM}};
  mem_37_MPORT_1_en_pipe_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  mem_37_MPORT_1_addr_pipe_0 = _RAND_113[3:0];
  _RAND_115 = {1{`RANDOM}};
  mem_38_MPORT_1_en_pipe_0 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  mem_38_MPORT_1_addr_pipe_0 = _RAND_116[3:0];
  _RAND_118 = {1{`RANDOM}};
  mem_39_MPORT_1_en_pipe_0 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  mem_39_MPORT_1_addr_pipe_0 = _RAND_119[3:0];
  _RAND_121 = {1{`RANDOM}};
  mem_40_MPORT_1_en_pipe_0 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  mem_40_MPORT_1_addr_pipe_0 = _RAND_122[3:0];
  _RAND_124 = {1{`RANDOM}};
  mem_41_MPORT_1_en_pipe_0 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  mem_41_MPORT_1_addr_pipe_0 = _RAND_125[3:0];
  _RAND_127 = {1{`RANDOM}};
  mem_42_MPORT_1_en_pipe_0 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  mem_42_MPORT_1_addr_pipe_0 = _RAND_128[3:0];
  _RAND_130 = {1{`RANDOM}};
  mem_43_MPORT_1_en_pipe_0 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  mem_43_MPORT_1_addr_pipe_0 = _RAND_131[3:0];
  _RAND_133 = {1{`RANDOM}};
  mem_44_MPORT_1_en_pipe_0 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  mem_44_MPORT_1_addr_pipe_0 = _RAND_134[3:0];
  _RAND_136 = {1{`RANDOM}};
  mem_45_MPORT_1_en_pipe_0 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  mem_45_MPORT_1_addr_pipe_0 = _RAND_137[3:0];
  _RAND_139 = {1{`RANDOM}};
  mem_46_MPORT_1_en_pipe_0 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  mem_46_MPORT_1_addr_pipe_0 = _RAND_140[3:0];
  _RAND_142 = {1{`RANDOM}};
  mem_47_MPORT_1_en_pipe_0 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  mem_47_MPORT_1_addr_pipe_0 = _RAND_143[3:0];
  _RAND_145 = {1{`RANDOM}};
  mem_48_MPORT_1_en_pipe_0 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  mem_48_MPORT_1_addr_pipe_0 = _RAND_146[3:0];
  _RAND_148 = {1{`RANDOM}};
  mem_49_MPORT_1_en_pipe_0 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  mem_49_MPORT_1_addr_pipe_0 = _RAND_149[3:0];
  _RAND_151 = {1{`RANDOM}};
  mem_50_MPORT_1_en_pipe_0 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  mem_50_MPORT_1_addr_pipe_0 = _RAND_152[3:0];
  _RAND_154 = {1{`RANDOM}};
  mem_51_MPORT_1_en_pipe_0 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  mem_51_MPORT_1_addr_pipe_0 = _RAND_155[3:0];
  _RAND_157 = {1{`RANDOM}};
  mem_52_MPORT_1_en_pipe_0 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  mem_52_MPORT_1_addr_pipe_0 = _RAND_158[3:0];
  _RAND_160 = {1{`RANDOM}};
  mem_53_MPORT_1_en_pipe_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  mem_53_MPORT_1_addr_pipe_0 = _RAND_161[3:0];
  _RAND_163 = {1{`RANDOM}};
  mem_54_MPORT_1_en_pipe_0 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  mem_54_MPORT_1_addr_pipe_0 = _RAND_164[3:0];
  _RAND_166 = {1{`RANDOM}};
  mem_55_MPORT_1_en_pipe_0 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  mem_55_MPORT_1_addr_pipe_0 = _RAND_167[3:0];
  _RAND_169 = {1{`RANDOM}};
  mem_56_MPORT_1_en_pipe_0 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  mem_56_MPORT_1_addr_pipe_0 = _RAND_170[3:0];
  _RAND_172 = {1{`RANDOM}};
  mem_57_MPORT_1_en_pipe_0 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  mem_57_MPORT_1_addr_pipe_0 = _RAND_173[3:0];
  _RAND_175 = {1{`RANDOM}};
  mem_58_MPORT_1_en_pipe_0 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  mem_58_MPORT_1_addr_pipe_0 = _RAND_176[3:0];
  _RAND_178 = {1{`RANDOM}};
  mem_59_MPORT_1_en_pipe_0 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  mem_59_MPORT_1_addr_pipe_0 = _RAND_179[3:0];
  _RAND_181 = {1{`RANDOM}};
  mem_60_MPORT_1_en_pipe_0 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  mem_60_MPORT_1_addr_pipe_0 = _RAND_182[3:0];
  _RAND_184 = {1{`RANDOM}};
  mem_61_MPORT_1_en_pipe_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  mem_61_MPORT_1_addr_pipe_0 = _RAND_185[3:0];
  _RAND_187 = {1{`RANDOM}};
  mem_62_MPORT_1_en_pipe_0 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  mem_62_MPORT_1_addr_pipe_0 = _RAND_188[3:0];
  _RAND_190 = {1{`RANDOM}};
  mem_63_MPORT_1_en_pipe_0 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  mem_63_MPORT_1_addr_pipe_0 = _RAND_191[3:0];
  _RAND_193 = {1{`RANDOM}};
  mem_64_MPORT_1_en_pipe_0 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  mem_64_MPORT_1_addr_pipe_0 = _RAND_194[3:0];
  _RAND_196 = {1{`RANDOM}};
  mem_65_MPORT_1_en_pipe_0 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  mem_65_MPORT_1_addr_pipe_0 = _RAND_197[3:0];
  _RAND_199 = {1{`RANDOM}};
  mem_66_MPORT_1_en_pipe_0 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  mem_66_MPORT_1_addr_pipe_0 = _RAND_200[3:0];
  _RAND_202 = {1{`RANDOM}};
  mem_67_MPORT_1_en_pipe_0 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  mem_67_MPORT_1_addr_pipe_0 = _RAND_203[3:0];
  _RAND_205 = {1{`RANDOM}};
  mem_68_MPORT_1_en_pipe_0 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  mem_68_MPORT_1_addr_pipe_0 = _RAND_206[3:0];
  _RAND_208 = {1{`RANDOM}};
  mem_69_MPORT_1_en_pipe_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  mem_69_MPORT_1_addr_pipe_0 = _RAND_209[3:0];
  _RAND_211 = {1{`RANDOM}};
  mem_70_MPORT_1_en_pipe_0 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  mem_70_MPORT_1_addr_pipe_0 = _RAND_212[3:0];
  _RAND_214 = {1{`RANDOM}};
  mem_71_MPORT_1_en_pipe_0 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  mem_71_MPORT_1_addr_pipe_0 = _RAND_215[3:0];
  _RAND_217 = {1{`RANDOM}};
  mem_72_MPORT_1_en_pipe_0 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  mem_72_MPORT_1_addr_pipe_0 = _RAND_218[3:0];
  _RAND_220 = {1{`RANDOM}};
  mem_73_MPORT_1_en_pipe_0 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  mem_73_MPORT_1_addr_pipe_0 = _RAND_221[3:0];
  _RAND_223 = {1{`RANDOM}};
  mem_74_MPORT_1_en_pipe_0 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  mem_74_MPORT_1_addr_pipe_0 = _RAND_224[3:0];
  _RAND_226 = {1{`RANDOM}};
  mem_75_MPORT_1_en_pipe_0 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  mem_75_MPORT_1_addr_pipe_0 = _RAND_227[3:0];
  _RAND_229 = {1{`RANDOM}};
  mem_76_MPORT_1_en_pipe_0 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  mem_76_MPORT_1_addr_pipe_0 = _RAND_230[3:0];
  _RAND_232 = {1{`RANDOM}};
  mem_77_MPORT_1_en_pipe_0 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  mem_77_MPORT_1_addr_pipe_0 = _RAND_233[3:0];
  _RAND_235 = {1{`RANDOM}};
  mem_78_MPORT_1_en_pipe_0 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  mem_78_MPORT_1_addr_pipe_0 = _RAND_236[3:0];
  _RAND_238 = {1{`RANDOM}};
  mem_79_MPORT_1_en_pipe_0 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  mem_79_MPORT_1_addr_pipe_0 = _RAND_239[3:0];
  _RAND_241 = {1{`RANDOM}};
  mem_80_MPORT_1_en_pipe_0 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  mem_80_MPORT_1_addr_pipe_0 = _RAND_242[3:0];
  _RAND_244 = {1{`RANDOM}};
  mem_81_MPORT_1_en_pipe_0 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  mem_81_MPORT_1_addr_pipe_0 = _RAND_245[3:0];
  _RAND_247 = {1{`RANDOM}};
  mem_82_MPORT_1_en_pipe_0 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  mem_82_MPORT_1_addr_pipe_0 = _RAND_248[3:0];
  _RAND_250 = {1{`RANDOM}};
  mem_83_MPORT_1_en_pipe_0 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  mem_83_MPORT_1_addr_pipe_0 = _RAND_251[3:0];
  _RAND_253 = {1{`RANDOM}};
  mem_84_MPORT_1_en_pipe_0 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  mem_84_MPORT_1_addr_pipe_0 = _RAND_254[3:0];
  _RAND_256 = {1{`RANDOM}};
  mem_85_MPORT_1_en_pipe_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  mem_85_MPORT_1_addr_pipe_0 = _RAND_257[3:0];
  _RAND_259 = {1{`RANDOM}};
  mem_86_MPORT_1_en_pipe_0 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  mem_86_MPORT_1_addr_pipe_0 = _RAND_260[3:0];
  _RAND_262 = {1{`RANDOM}};
  mem_87_MPORT_1_en_pipe_0 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  mem_87_MPORT_1_addr_pipe_0 = _RAND_263[3:0];
  _RAND_265 = {1{`RANDOM}};
  mem_88_MPORT_1_en_pipe_0 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  mem_88_MPORT_1_addr_pipe_0 = _RAND_266[3:0];
  _RAND_268 = {1{`RANDOM}};
  mem_89_MPORT_1_en_pipe_0 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  mem_89_MPORT_1_addr_pipe_0 = _RAND_269[3:0];
  _RAND_271 = {1{`RANDOM}};
  mem_90_MPORT_1_en_pipe_0 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  mem_90_MPORT_1_addr_pipe_0 = _RAND_272[3:0];
  _RAND_274 = {1{`RANDOM}};
  mem_91_MPORT_1_en_pipe_0 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  mem_91_MPORT_1_addr_pipe_0 = _RAND_275[3:0];
  _RAND_277 = {1{`RANDOM}};
  mem_92_MPORT_1_en_pipe_0 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  mem_92_MPORT_1_addr_pipe_0 = _RAND_278[3:0];
  _RAND_280 = {1{`RANDOM}};
  mem_93_MPORT_1_en_pipe_0 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  mem_93_MPORT_1_addr_pipe_0 = _RAND_281[3:0];
  _RAND_283 = {1{`RANDOM}};
  mem_94_MPORT_1_en_pipe_0 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  mem_94_MPORT_1_addr_pipe_0 = _RAND_284[3:0];
  _RAND_286 = {1{`RANDOM}};
  mem_95_MPORT_1_en_pipe_0 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  mem_95_MPORT_1_addr_pipe_0 = _RAND_287[3:0];
  _RAND_289 = {1{`RANDOM}};
  mem_96_MPORT_1_en_pipe_0 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  mem_96_MPORT_1_addr_pipe_0 = _RAND_290[3:0];
  _RAND_292 = {1{`RANDOM}};
  mem_97_MPORT_1_en_pipe_0 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  mem_97_MPORT_1_addr_pipe_0 = _RAND_293[3:0];
  _RAND_295 = {1{`RANDOM}};
  mem_98_MPORT_1_en_pipe_0 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  mem_98_MPORT_1_addr_pipe_0 = _RAND_296[3:0];
  _RAND_298 = {1{`RANDOM}};
  mem_99_MPORT_1_en_pipe_0 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  mem_99_MPORT_1_addr_pipe_0 = _RAND_299[3:0];
  _RAND_301 = {1{`RANDOM}};
  mem_100_MPORT_1_en_pipe_0 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  mem_100_MPORT_1_addr_pipe_0 = _RAND_302[3:0];
  _RAND_304 = {1{`RANDOM}};
  mem_101_MPORT_1_en_pipe_0 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  mem_101_MPORT_1_addr_pipe_0 = _RAND_305[3:0];
  _RAND_307 = {1{`RANDOM}};
  mem_102_MPORT_1_en_pipe_0 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  mem_102_MPORT_1_addr_pipe_0 = _RAND_308[3:0];
  _RAND_310 = {1{`RANDOM}};
  mem_103_MPORT_1_en_pipe_0 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  mem_103_MPORT_1_addr_pipe_0 = _RAND_311[3:0];
  _RAND_313 = {1{`RANDOM}};
  mem_104_MPORT_1_en_pipe_0 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  mem_104_MPORT_1_addr_pipe_0 = _RAND_314[3:0];
  _RAND_316 = {1{`RANDOM}};
  mem_105_MPORT_1_en_pipe_0 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  mem_105_MPORT_1_addr_pipe_0 = _RAND_317[3:0];
  _RAND_319 = {1{`RANDOM}};
  mem_106_MPORT_1_en_pipe_0 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  mem_106_MPORT_1_addr_pipe_0 = _RAND_320[3:0];
  _RAND_322 = {1{`RANDOM}};
  mem_107_MPORT_1_en_pipe_0 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  mem_107_MPORT_1_addr_pipe_0 = _RAND_323[3:0];
  _RAND_325 = {1{`RANDOM}};
  mem_108_MPORT_1_en_pipe_0 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  mem_108_MPORT_1_addr_pipe_0 = _RAND_326[3:0];
  _RAND_328 = {1{`RANDOM}};
  mem_109_MPORT_1_en_pipe_0 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  mem_109_MPORT_1_addr_pipe_0 = _RAND_329[3:0];
  _RAND_331 = {1{`RANDOM}};
  mem_110_MPORT_1_en_pipe_0 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  mem_110_MPORT_1_addr_pipe_0 = _RAND_332[3:0];
  _RAND_334 = {1{`RANDOM}};
  mem_111_MPORT_1_en_pipe_0 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  mem_111_MPORT_1_addr_pipe_0 = _RAND_335[3:0];
  _RAND_337 = {1{`RANDOM}};
  mem_112_MPORT_1_en_pipe_0 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  mem_112_MPORT_1_addr_pipe_0 = _RAND_338[3:0];
  _RAND_340 = {1{`RANDOM}};
  mem_113_MPORT_1_en_pipe_0 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  mem_113_MPORT_1_addr_pipe_0 = _RAND_341[3:0];
  _RAND_343 = {1{`RANDOM}};
  mem_114_MPORT_1_en_pipe_0 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  mem_114_MPORT_1_addr_pipe_0 = _RAND_344[3:0];
  _RAND_346 = {1{`RANDOM}};
  mem_115_MPORT_1_en_pipe_0 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  mem_115_MPORT_1_addr_pipe_0 = _RAND_347[3:0];
  _RAND_349 = {1{`RANDOM}};
  mem_116_MPORT_1_en_pipe_0 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  mem_116_MPORT_1_addr_pipe_0 = _RAND_350[3:0];
  _RAND_352 = {1{`RANDOM}};
  mem_117_MPORT_1_en_pipe_0 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  mem_117_MPORT_1_addr_pipe_0 = _RAND_353[3:0];
  _RAND_355 = {1{`RANDOM}};
  mem_118_MPORT_1_en_pipe_0 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  mem_118_MPORT_1_addr_pipe_0 = _RAND_356[3:0];
  _RAND_358 = {1{`RANDOM}};
  mem_119_MPORT_1_en_pipe_0 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  mem_119_MPORT_1_addr_pipe_0 = _RAND_359[3:0];
  _RAND_361 = {1{`RANDOM}};
  mem_120_MPORT_1_en_pipe_0 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  mem_120_MPORT_1_addr_pipe_0 = _RAND_362[3:0];
  _RAND_364 = {1{`RANDOM}};
  mem_121_MPORT_1_en_pipe_0 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  mem_121_MPORT_1_addr_pipe_0 = _RAND_365[3:0];
  _RAND_367 = {1{`RANDOM}};
  mem_122_MPORT_1_en_pipe_0 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  mem_122_MPORT_1_addr_pipe_0 = _RAND_368[3:0];
  _RAND_370 = {1{`RANDOM}};
  mem_123_MPORT_1_en_pipe_0 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  mem_123_MPORT_1_addr_pipe_0 = _RAND_371[3:0];
  _RAND_373 = {1{`RANDOM}};
  mem_124_MPORT_1_en_pipe_0 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  mem_124_MPORT_1_addr_pipe_0 = _RAND_374[3:0];
  _RAND_376 = {1{`RANDOM}};
  mem_125_MPORT_1_en_pipe_0 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  mem_125_MPORT_1_addr_pipe_0 = _RAND_377[3:0];
  _RAND_379 = {1{`RANDOM}};
  mem_126_MPORT_1_en_pipe_0 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  mem_126_MPORT_1_addr_pipe_0 = _RAND_380[3:0];
  _RAND_382 = {1{`RANDOM}};
  mem_127_MPORT_1_en_pipe_0 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  mem_127_MPORT_1_addr_pipe_0 = _RAND_383[3:0];
  _RAND_384 = {1{`RANDOM}};
  counter = _RAND_384[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
