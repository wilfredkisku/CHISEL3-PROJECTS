module FP16Add(
  input         clock,
  input         reset,
  input  [15:0] io_a,
  input  [15:0] io_b,
  output [15:0] io_result
);
  wire  signA = io_a[15]; // @[FP16Add.scala 13:18]
  wire [4:0] expA = io_a[14:10]; // @[FP16Add.scala 14:22]
  wire [9:0] sigA = io_a[9:0]; // @[FP16Add.scala 15:25]
  wire  signB = io_b[15]; // @[FP16Add.scala 13:18]
  wire [4:0] expB = io_b[14:10]; // @[FP16Add.scala 14:22]
  wire [9:0] sigB = io_b[9:0]; // @[FP16Add.scala 15:25]
  wire  _zeroFlagA_T = expA == 5'h0; // @[FP16Add.scala 38:24]
  wire  _zeroFlagA_T_1 = sigA == 10'h0; // @[FP16Add.scala 38:40]
  wire  zeroFlagA = expA == 5'h0 & sigA == 10'h0; // @[FP16Add.scala 38:32]
  wire  _zeroFlagB_T = expB == 5'h0; // @[FP16Add.scala 39:24]
  wire  _zeroFlagB_T_1 = sigB == 10'h0; // @[FP16Add.scala 39:40]
  wire  zeroFlagB = expB == 5'h0 & sigB == 10'h0; // @[FP16Add.scala 39:32]
  wire  infFlagA = expA == 5'h1f & _zeroFlagA_T_1; // @[FP16Add.scala 44:38]
  wire  infFlagB = expB == 5'h1f & _zeroFlagB_T_1; // @[FP16Add.scala 45:38]
  wire  subNormA = _zeroFlagA_T & sigA != 10'h0; // @[FP16Add.scala 47:31]
  wire  subNormB = _zeroFlagB_T & sigB != 10'h0; // @[FP16Add.scala 48:31]
  wire [15:0] _io_result_T = infFlagA ? io_a : io_b; // @[FP16Add.scala 73:25]
  wire [15:0] _GEN_0 = infFlagA & infFlagB & signA != signB ? 16'h7fff : _io_result_T; // @[FP16Add.scala 67:54 69:19 73:19]
  wire [9:0] _GEN_18 = {{5'd0}, expA}; // @[FP16Add.scala 75:49]
  wire [9:0] _GEN_19 = {{5'd0}, expB}; // @[FP16Add.scala 75:106]
  wire  _T_20 = ~signA; // @[FP16Add.scala 86:22]
  wire  _T_21 = ~signB; // @[FP16Add.scala 86:39]
  wire [10:0] _io_result_T_1 = {1'h1,sigA}; // @[Cat.scala 33:92]
  wire [10:0] _io_result_T_2 = {1'h1,sigB}; // @[Cat.scala 33:92]
  wire [11:0] _io_result_T_3 = _io_result_T_1 + _io_result_T_2; // @[FP16Add.scala 89:46]
  wire [4:0] _io_result_T_7 = expA + 5'h1; // @[FP16Add.scala 89:94]
  wire [15:0] _io_result_T_12 = {signA,_io_result_T_7,_io_result_T_3[10:1]}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_17 = {signA,expA,_io_result_T_3[9:0]}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_18 = _io_result_T_3[11] ? _io_result_T_12 : _io_result_T_17; // @[FP16Add.scala 89:29]
  wire  _io_result_T_19 = sigB >= sigA; // @[FP16Add.scala 92:35]
  wire [10:0] _io_result_T_23 = _io_result_T_2 - _io_result_T_1; // @[FP16Add.scala 92:75]
  wire [15:0] _io_result_T_25 = {1'h0,expB,_io_result_T_23[9:0]}; // @[Cat.scala 33:92]
  wire [10:0] _io_result_T_29 = _io_result_T_1 - _io_result_T_2; // @[FP16Add.scala 92:131]
  wire [15:0] _io_result_T_31 = {1'h1,expA,_io_result_T_29[9:0]}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_32 = sigB >= sigA ? _io_result_T_25 : _io_result_T_31; // @[FP16Add.scala 92:29]
  wire [15:0] _io_result_T_39 = {1'h1,expB,_io_result_T_23[9:0]}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_45 = {1'h0,expA,_io_result_T_29[9:0]}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_46 = _io_result_T_19 ? _io_result_T_39 : _io_result_T_45; // @[FP16Add.scala 94:29]
  wire [15:0] _GEN_1 = _T_20 & signB ? _io_result_T_46 : _io_result_T_18; // @[FP16Add.scala 93:53 94:23 96:23]
  wire [15:0] _GEN_2 = signA & _T_21 ? _io_result_T_32 : _GEN_1; // @[FP16Add.scala 90:53 92:23]
  wire [15:0] _GEN_3 = ~signA & ~signB ? _io_result_T_18 : _GEN_2; // @[FP16Add.scala 86:47 89:23]
  wire [4:0] _io_result_T_68 = expA - expB; // @[FP16Add.scala 106:107]
  wire [9:0] _io_result_T_69 = sigB >> _io_result_T_68; // @[FP16Add.scala 106:99]
  wire [10:0] _io_result_T_70 = {1'h0,_io_result_T_69}; // @[Cat.scala 33:92]
  wire [10:0] _io_result_T_72 = _io_result_T_1 + _io_result_T_70; // @[FP16Add.scala 106:83]
  wire [16:0] _io_result_T_73 = {1'h0,expA,_io_result_T_72}; // @[Cat.scala 33:92]
  wire [10:0] _io_result_T_78 = {1'h1,_io_result_T_69}; // @[Cat.scala 33:92]
  wire [10:0] _io_result_T_80 = _io_result_T_1 - _io_result_T_78; // @[FP16Add.scala 106:147]
  wire [16:0] _io_result_T_81 = {1'h0,expA,_io_result_T_80}; // @[Cat.scala 33:92]
  wire [16:0] _io_result_T_82 = _T_21 ? _io_result_T_73 : _io_result_T_81; // @[FP16Add.scala 106:37]
  wire [10:0] _io_result_T_90 = _io_result_T_1 - _io_result_T_70; // @[FP16Add.scala 108:79]
  wire [16:0] _io_result_T_91 = {1'h1,expA,_io_result_T_90}; // @[Cat.scala 33:92]
  wire [10:0] _io_result_T_98 = _io_result_T_1 + _io_result_T_78; // @[FP16Add.scala 108:143]
  wire [16:0] _io_result_T_99 = {1'h1,expA,_io_result_T_98}; // @[Cat.scala 33:92]
  wire [16:0] _io_result_T_100 = _T_21 ? _io_result_T_91 : _io_result_T_99; // @[FP16Add.scala 108:33]
  wire [16:0] _GEN_4 = _T_20 ? _io_result_T_82 : _io_result_T_100; // @[FP16Add.scala 105:34 106:31 108:27]
  wire [4:0] _io_result_T_104 = expB - expA; // @[FP16Add.scala 114:99]
  wire [9:0] _io_result_T_105 = sigA >> _io_result_T_104; // @[FP16Add.scala 114:91]
  wire [10:0] _io_result_T_106 = {1'h0,_io_result_T_105}; // @[Cat.scala 33:92]
  wire [10:0] _io_result_T_108 = _io_result_T_2 + _io_result_T_106; // @[FP16Add.scala 114:75]
  wire [16:0] _io_result_T_109 = {1'h0,expB,_io_result_T_108}; // @[Cat.scala 33:92]
  wire [10:0] _io_result_T_114 = {1'h1,_io_result_T_105}; // @[Cat.scala 33:92]
  wire [10:0] _io_result_T_116 = _io_result_T_2 - _io_result_T_114; // @[FP16Add.scala 114:139]
  wire [16:0] _io_result_T_117 = {1'h0,expB,_io_result_T_116}; // @[Cat.scala 33:92]
  wire [16:0] _io_result_T_118 = _T_20 ? _io_result_T_109 : _io_result_T_117; // @[FP16Add.scala 114:29]
  wire [10:0] _io_result_T_126 = _io_result_T_2 - _io_result_T_106; // @[FP16Add.scala 116:75]
  wire [16:0] _io_result_T_127 = {1'h1,expB,_io_result_T_126}; // @[Cat.scala 33:92]
  wire [10:0] _io_result_T_134 = _io_result_T_2 + _io_result_T_114; // @[FP16Add.scala 116:139]
  wire [16:0] _io_result_T_135 = {1'h1,expB,_io_result_T_134}; // @[Cat.scala 33:92]
  wire [16:0] _io_result_T_136 = _T_20 ? _io_result_T_127 : _io_result_T_135; // @[FP16Add.scala 116:29]
  wire [16:0] _GEN_5 = _T_21 ? _io_result_T_118 : _io_result_T_136; // @[FP16Add.scala 113:30 114:23 116:23]
  wire [16:0] _GEN_6 = expA > expB ? _GEN_4 : _GEN_5; // @[FP16Add.scala 98:33]
  wire [16:0] _GEN_7 = expA == expB ? {{1'd0}, _GEN_3} : _GEN_6; // @[FP16Add.scala 83:29]
  wire [10:0] _io_result_T_138 = {1'h0,sigB}; // @[Cat.scala 33:92]
  wire [10:0] _io_result_T_139 = {1'h0,sigA}; // @[Cat.scala 33:92]
  wire [10:0] _io_result_T_141 = _io_result_T_138 + _io_result_T_139; // @[FP16Add.scala 125:75]
  wire [16:0] _io_result_T_142 = {1'h1,expB,_io_result_T_141}; // @[Cat.scala 33:92]
  wire [10:0] _io_result_T_146 = _io_result_T_138 - _io_result_T_139; // @[FP16Add.scala 125:124]
  wire [16:0] _io_result_T_147 = {1'h1,expB,_io_result_T_146}; // @[Cat.scala 33:92]
  wire [16:0] _io_result_T_148 = signA ? _io_result_T_142 : _io_result_T_147; // @[FP16Add.scala 125:29]
  wire [16:0] _io_result_T_154 = {1'h0,expB,_io_result_T_146}; // @[Cat.scala 33:92]
  wire [16:0] _io_result_T_159 = {1'h0,expB,_io_result_T_141}; // @[Cat.scala 33:92]
  wire [16:0] _io_result_T_160 = signA ? _io_result_T_154 : _io_result_T_159; // @[FP16Add.scala 128:31]
  wire [16:0] _GEN_8 = signB ? _io_result_T_148 : _io_result_T_160; // @[FP16Add.scala 124:30 125:23 128:25]
  wire [10:0] _io_result_T_165 = _io_result_T_139 + _io_result_T_138; // @[FP16Add.scala 133:75]
  wire [16:0] _io_result_T_166 = {1'h1,expA,_io_result_T_165}; // @[Cat.scala 33:92]
  wire [10:0] _io_result_T_170 = _io_result_T_139 - _io_result_T_138; // @[FP16Add.scala 133:124]
  wire [16:0] _io_result_T_171 = {1'h1,expA,_io_result_T_170}; // @[Cat.scala 33:92]
  wire [16:0] _io_result_T_172 = signB ? _io_result_T_166 : _io_result_T_171; // @[FP16Add.scala 133:29]
  wire [16:0] _io_result_T_178 = {1'h0,expA,_io_result_T_170}; // @[Cat.scala 33:92]
  wire [16:0] _io_result_T_183 = {1'h0,expA,_io_result_T_165}; // @[Cat.scala 33:92]
  wire [16:0] _io_result_T_184 = signB ? _io_result_T_178 : _io_result_T_183; // @[FP16Add.scala 136:31]
  wire [16:0] _GEN_9 = signA ? _io_result_T_172 : _io_result_T_184; // @[FP16Add.scala 132:30 133:23 136:25]
  wire [16:0] _GEN_10 = sigA < sigB ? _GEN_8 : _GEN_9; // @[FP16Add.scala 123:26]
  wire [16:0] _GEN_11 = subNormA & subNormB ? _GEN_10 : 17'h0; // @[FP16Add.scala 121:38 142:19]
  wire [16:0] _GEN_12 = ~subNormA & ~subNormB ? _GEN_7 : _GEN_11; // @[FP16Add.scala 80:34]
  wire [16:0] _GEN_13 = sigA == 10'h1f & _GEN_18 == 10'h3ff | sigB == 10'h1f & _GEN_19 == 10'h3ff ? 17'h7fff : _GEN_12; // @[FP16Add.scala 75:128 76:17]
  wire [16:0] _GEN_14 = infFlagA | infFlagB ? {{1'd0}, _GEN_0} : _GEN_13; // @[FP16Add.scala 65:38]
  wire [16:0] _GEN_15 = zeroFlagA & ~zeroFlagB ? {{1'd0}, io_b} : _GEN_14; // @[FP16Add.scala 62:41 64:17]
  wire [16:0] _GEN_16 = ~zeroFlagA & zeroFlagB ? {{1'd0}, io_a} : _GEN_15; // @[FP16Add.scala 59:40 61:17]
  wire [16:0] _GEN_17 = zeroFlagA & zeroFlagB ? 17'h0 : _GEN_16; // @[FP16Add.scala 55:32 57:17]
  assign io_result = _GEN_17[15:0];
endmodule
