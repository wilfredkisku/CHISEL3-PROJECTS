module FP8_ADD(
  input        clock,
  input        reset,
  input  [7:0] io_inputA,
  input  [7:0] io_inputB,
  output [7:0] io_output
);
  wire  signA = io_inputA[7]; // @[FP8_ADD.scala 13:18]
  wire [4:0] expA = io_inputA[6:2]; // @[FP8_ADD.scala 14:22]
  wire [1:0] sigA = io_inputA[1:0]; // @[FP8_ADD.scala 15:25]
  wire  signB = io_inputB[7]; // @[FP8_ADD.scala 13:18]
  wire [4:0] expB = io_inputB[6:2]; // @[FP8_ADD.scala 14:22]
  wire [1:0] sigB = io_inputB[1:0]; // @[FP8_ADD.scala 15:25]
  wire  _infFlagA_T = expA == 5'h1f; // @[FP8_ADD.scala 24:23]
  wire  _infFlagA_T_1 = sigA == 2'h0; // @[FP8_ADD.scala 24:46]
  wire  infFlagA = expA == 5'h1f & sigA == 2'h0; // @[FP8_ADD.scala 24:38]
  wire  _infFlagB_T = expB == 5'h1f; // @[FP8_ADD.scala 25:23]
  wire  _infFlagB_T_1 = sigB == 2'h0; // @[FP8_ADD.scala 25:46]
  wire  infFlagB = expB == 5'h1f & sigB == 2'h0; // @[FP8_ADD.scala 25:38]
  wire  _zeroFlagA_T = expA == 5'h0; // @[FP8_ADD.scala 28:24]
  wire  zeroFlagA = expA == 5'h0 & _infFlagA_T_1; // @[FP8_ADD.scala 28:39]
  wire  _zeroFlagB_T = expB == 5'h0; // @[FP8_ADD.scala 29:24]
  wire  zeroFlagB = expB == 5'h0 & _infFlagB_T_1; // @[FP8_ADD.scala 29:39]
  wire  _nanFlagA_T_1 = sigA != 2'h0; // @[FP8_ADD.scala 32:46]
  wire  nanFlagA = _infFlagA_T & sigA != 2'h0; // @[FP8_ADD.scala 32:38]
  wire  _nanFlagB_T_1 = sigB != 2'h0; // @[FP8_ADD.scala 33:46]
  wire  nanFlagB = _infFlagB_T & sigB != 2'h0; // @[FP8_ADD.scala 33:38]
  wire  subFlagA = _zeroFlagA_T & _nanFlagA_T_1; // @[FP8_ADD.scala 36:38]
  wire  subFlagB = _zeroFlagB_T & _nanFlagB_T_1; // @[FP8_ADD.scala 37:38]
  wire [7:0] _io_output_T = infFlagA ? io_inputA : io_inputB; // @[FP8_ADD.scala 55:23]
  wire [7:0] _GEN_0 = infFlagA & infFlagB & signA != signB ? 8'h7f : _io_output_T; // @[FP8_ADD.scala 52:53 53:17 55:17]
  wire [2:0] _ovrChk_a_T = {1'h1,sigA}; // @[Cat.scala 33:92]
  wire [2:0] _ovrChk_a_T_1 = {1'h1,sigB}; // @[Cat.scala 33:92]
  wire [4:0] _ovrChk_a_T_3 = expA - expB; // @[FP8_ADD.scala 80:64]
  wire [2:0] _ovrChk_a_T_4 = _ovrChk_a_T_1 >> _ovrChk_a_T_3; // @[FP8_ADD.scala 80:55]
  wire [3:0] _ovrChk_a_T_5 = _ovrChk_a_T + _ovrChk_a_T_4; // @[FP8_ADD.scala 80:36]
  wire [2:0] _ovrChk_s_T_6 = _ovrChk_a_T - _ovrChk_a_T_4; // @[FP8_ADD.scala 81:36]
  wire  _io_output_T_1 = ~signA; // @[FP8_ADD.scala 82:32]
  wire  _io_output_T_2 = ~signB; // @[FP8_ADD.scala 82:68]
  wire [4:0] _ovrChk_a_T_9 = expB - expA; // @[FP8_ADD.scala 85:64]
  wire [2:0] _ovrChk_a_T_10 = _ovrChk_a_T >> _ovrChk_a_T_9; // @[FP8_ADD.scala 85:55]
  wire [3:0] _ovrChk_a_T_11 = _ovrChk_a_T_1 + _ovrChk_a_T_10; // @[FP8_ADD.scala 85:36]
  wire [3:0] _GEN_1 = expA > expB ? _ovrChk_a_T_5 : _ovrChk_a_T_11; // @[FP8_ADD.scala 78:24 80:18 85:18]
  wire [3:0] _GEN_4 = ~subFlagA & ~subFlagB ? _GEN_1 : 4'h0; // @[FP8_ADD.scala 43:12 69:39]
  wire [3:0] _GEN_8 = subFlagA & subFlagB ? 4'h0 : _GEN_4; // @[FP8_ADD.scala 43:12 61:31]
  wire [3:0] _GEN_11 = nanFlagA | nanFlagB ? 4'h0 : _GEN_8; // @[FP8_ADD.scala 43:12 57:35]
  wire [3:0] _GEN_14 = infFlagA | infFlagB ? 4'h0 : _GEN_11; // @[FP8_ADD.scala 43:12 50:35]
  wire [3:0] ovrChk_a = zeroFlagA & zeroFlagB ? 4'h0 : _GEN_14; // @[FP8_ADD.scala 43:12 47:32]
  wire [2:0] _ovrChk_s_T_13 = _ovrChk_a_T_1 - _ovrChk_a_T_10; // @[FP8_ADD.scala 86:36]
  wire [2:0] _GEN_2 = expA > expB ? _ovrChk_s_T_6 : _ovrChk_s_T_13; // @[FP8_ADD.scala 78:24 81:18 86:18]
  wire [2:0] _GEN_5 = ~subFlagA & ~subFlagB ? _GEN_2 : 3'h0; // @[FP8_ADD.scala 44:12 69:39]
  wire [2:0] _GEN_9 = subFlagA & subFlagB ? 3'h0 : _GEN_5; // @[FP8_ADD.scala 44:12 61:31]
  wire [2:0] _GEN_12 = nanFlagA | nanFlagB ? 3'h0 : _GEN_9; // @[FP8_ADD.scala 44:12 57:35]
  wire [2:0] _GEN_15 = infFlagA | infFlagB ? 3'h0 : _GEN_12; // @[FP8_ADD.scala 44:12 50:35]
  wire [2:0] _GEN_18 = zeroFlagA & zeroFlagB ? 3'h0 : _GEN_15; // @[FP8_ADD.scala 44:12 47:32]
  wire [3:0] ovrChk_s = {{1'd0}, _GEN_18}; // @[FP8_ADD.scala 41:22]
  wire [1:0] _io_output_T_5 = ~signB ? ovrChk_a[1:0] : ovrChk_s[1:0]; // @[FP8_ADD.scala 82:61]
  wire [7:0] _io_output_T_6 = {signA,expA,_io_output_T_5}; // @[Cat.scala 33:92]
  wire [1:0] _io_output_T_10 = ~signB ? ovrChk_s[1:0] : ovrChk_a[1:0]; // @[FP8_ADD.scala 82:129]
  wire [7:0] _io_output_T_11 = {signA,expA,_io_output_T_10}; // @[Cat.scala 33:92]
  wire [7:0] _io_output_T_12 = ~signA ? _io_output_T_6 : _io_output_T_11; // @[FP8_ADD.scala 82:25]
  wire [1:0] _io_output_T_17 = _io_output_T_1 ? ovrChk_a[1:0] : ovrChk_s[1:0]; // @[FP8_ADD.scala 87:61]
  wire [7:0] _io_output_T_18 = {signB,expB,_io_output_T_17}; // @[Cat.scala 33:92]
  wire [1:0] _io_output_T_22 = _io_output_T_1 ? ovrChk_s[1:0] : ovrChk_a[1:0]; // @[FP8_ADD.scala 87:129]
  wire [7:0] _io_output_T_23 = {signB,expB,_io_output_T_22}; // @[Cat.scala 33:92]
  wire [7:0] _io_output_T_24 = _io_output_T_2 ? _io_output_T_18 : _io_output_T_23; // @[FP8_ADD.scala 87:25]
  wire [7:0] _GEN_3 = expA > expB ? _io_output_T_12 : _io_output_T_24; // @[FP8_ADD.scala 78:24 82:19 87:19]
  wire [7:0] _GEN_6 = ~subFlagA & ~subFlagB ? _GEN_3 : 8'h0; // @[FP8_ADD.scala 69:39 96:17]
  wire [7:0] _GEN_7 = subFlagA & subFlagB ? 8'h0 : _GEN_6; // @[FP8_ADD.scala 61:31 65:17]
  wire [7:0] _GEN_10 = nanFlagA | nanFlagB ? 8'h7f : _GEN_7; // @[FP8_ADD.scala 57:35 58:15]
  wire [7:0] _GEN_13 = infFlagA | infFlagB ? _GEN_0 : _GEN_10; // @[FP8_ADD.scala 50:35]
  assign io_output = zeroFlagA & zeroFlagB ? 8'h0 : _GEN_13; // @[FP8_ADD.scala 47:32 49:15]
endmodule
