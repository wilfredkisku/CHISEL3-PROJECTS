module FP16Add(
  input         clock,
  input         reset,
  input  [15:0] io_a,
  input  [15:0] io_b,
  output [15:0] io_result
);
  wire  signA = io_a[15]; // @[FP16Add.scala 13:18]
  wire [4:0] expA = io_a[14:10]; // @[FP16Add.scala 14:22]
  wire [9:0] sigA = io_a[9:0]; // @[FP16Add.scala 15:25]
  wire  signB = io_b[15]; // @[FP16Add.scala 13:18]
  wire [4:0] expB = io_b[14:10]; // @[FP16Add.scala 14:22]
  wire [9:0] sigB = io_b[9:0]; // @[FP16Add.scala 15:25]
  wire  _zeroFlagA_T_1 = sigA == 10'h0; // @[FP16Add.scala 38:40]
  wire  zeroFlagA = expA == 5'h0 & sigA == 10'h0; // @[FP16Add.scala 38:32]
  wire  _zeroFlagB_T_1 = sigB == 10'h0; // @[FP16Add.scala 39:40]
  wire  zeroFlagB = expB == 5'h0 & sigB == 10'h0; // @[FP16Add.scala 39:32]
  wire  infFlagA = expA == 5'h1f & _zeroFlagA_T_1; // @[FP16Add.scala 41:38]
  wire  infFlagB = expB == 5'h1f & _zeroFlagB_T_1; // @[FP16Add.scala 42:38]
  wire [15:0] _io_result_T = infFlagA ? io_a : io_b; // @[FP16Add.scala 64:25]
  wire [15:0] _GEN_0 = infFlagA & infFlagB & signA != signB ? 16'h7fff : _io_result_T; // @[FP16Add.scala 58:54 60:19 64:19]
  wire [10:0] _norm_T = {1'h1,sigB}; // @[Cat.scala 33:92]
  wire [4:0] _norm_T_2 = expA - expB; // @[FP16Add.scala 71:44]
  wire [10:0] _norm_T_3 = _norm_T >> _norm_T_2; // @[FP16Add.scala 71:35]
  wire  _io_result_T_1 = ~signA; // @[FP16Add.scala 72:32]
  wire  _io_result_T_2 = ~signB; // @[FP16Add.scala 72:51]
  wire [10:0] _norm_T_5 = {1'h1,sigA}; // @[Cat.scala 33:92]
  wire [4:0] _norm_T_7 = expB - expA; // @[FP16Add.scala 86:44]
  wire [10:0] _norm_T_8 = _norm_T_5 >> _norm_T_7; // @[FP16Add.scala 86:35]
  wire [9:0] _GEN_4 = expA == expB ? 10'h0 : _norm_T_8[10:1]; // @[FP16Add.scala 73:32 45:8 86:14]
  wire [9:0] _GEN_5 = expA > expB ? _norm_T_3[10:1] : _GEN_4; // @[FP16Add.scala 69:24 71:14]
  wire [9:0] _GEN_8 = infFlagA | infFlagB ? 10'h0 : _GEN_5; // @[FP16Add.scala 56:38 45:8]
  wire [9:0] _GEN_10 = zeroFlagA & ~zeroFlagB ? 10'h0 : _GEN_8; // @[FP16Add.scala 53:41 45:8]
  wire [9:0] _GEN_12 = ~zeroFlagA & zeroFlagB ? 10'h0 : _GEN_10; // @[FP16Add.scala 50:40 45:8]
  wire [9:0] norm = zeroFlagA & zeroFlagB ? 10'h0 : _GEN_12; // @[FP16Add.scala 46:32 45:8]
  wire [9:0] _io_result_T_4 = sigA + norm; // @[FP16Add.scala 72:78]
  wire [15:0] _io_result_T_5 = {1'h0,expA,_io_result_T_4}; // @[Cat.scala 33:92]
  wire [9:0] _io_result_T_7 = sigA - norm; // @[FP16Add.scala 72:107]
  wire [15:0] _io_result_T_8 = {1'h0,expA,_io_result_T_7}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_9 = ~signB ? _io_result_T_5 : _io_result_T_8; // @[FP16Add.scala 72:44]
  wire [15:0] _io_result_T_13 = {1'h1,expA,_io_result_T_7}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_16 = {1'h1,expA,_io_result_T_4}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_17 = ~signB ? _io_result_T_13 : _io_result_T_16; // @[FP16Add.scala 72:120]
  wire [15:0] _io_result_T_18 = ~signA ? _io_result_T_9 : _io_result_T_17; // @[FP16Add.scala 72:25]
  wire [9:0] _io_result_T_22 = sigA + sigB; // @[FP16Add.scala 76:80]
  wire [15:0] _io_result_T_23 = {1'h0,expA,_io_result_T_22}; // @[Cat.scala 33:92]
  wire [9:0] _io_result_T_25 = sigA - sigB; // @[FP16Add.scala 76:109]
  wire [15:0] _io_result_T_26 = {1'h0,expA,_io_result_T_25}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_27 = _io_result_T_2 ? _io_result_T_23 : _io_result_T_26; // @[FP16Add.scala 76:46]
  wire [15:0] _io_result_T_31 = {1'h1,expA,_io_result_T_25}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_34 = {1'h1,expA,_io_result_T_22}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_35 = _io_result_T_2 ? _io_result_T_31 : _io_result_T_34; // @[FP16Add.scala 76:122]
  wire [15:0] _io_result_T_36 = _io_result_T_1 ? _io_result_T_27 : _io_result_T_35; // @[FP16Add.scala 76:27]
  wire [9:0] _io_result_T_40 = sigB + sigA; // @[FP16Add.scala 79:82]
  wire [15:0] _io_result_T_41 = {1'h0,expB,_io_result_T_40}; // @[Cat.scala 33:92]
  wire [9:0] _io_result_T_43 = sigB - sigA; // @[FP16Add.scala 79:111]
  wire [15:0] _io_result_T_44 = {1'h0,expB,_io_result_T_43}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_45 = _io_result_T_1 ? _io_result_T_41 : _io_result_T_44; // @[FP16Add.scala 79:48]
  wire [15:0] _io_result_T_49 = {1'h1,expB,_io_result_T_43}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_52 = {1'h1,expB,_io_result_T_40}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_53 = _io_result_T_1 ? _io_result_T_49 : _io_result_T_52; // @[FP16Add.scala 79:124]
  wire [15:0] _io_result_T_54 = _io_result_T_2 ? _io_result_T_45 : _io_result_T_53; // @[FP16Add.scala 79:29]
  wire [15:0] _GEN_1 = sigB > sigA ? _io_result_T_54 : 16'h0; // @[FP16Add.scala 78:34 79:23 82:22]
  wire [15:0] _GEN_2 = sigA > sigB ? _io_result_T_36 : _GEN_1; // @[FP16Add.scala 75:28 76:21]
  wire [9:0] _io_result_T_58 = sigB + norm; // @[FP16Add.scala 87:78]
  wire [15:0] _io_result_T_59 = {1'h0,expB,_io_result_T_58}; // @[Cat.scala 33:92]
  wire [9:0] _io_result_T_61 = sigB - norm; // @[FP16Add.scala 87:107]
  wire [15:0] _io_result_T_62 = {1'h0,expB,_io_result_T_61}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_63 = _io_result_T_1 ? _io_result_T_59 : _io_result_T_62; // @[FP16Add.scala 87:44]
  wire [15:0] _io_result_T_67 = {1'h1,expB,_io_result_T_61}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_70 = {1'h1,expB,_io_result_T_58}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_71 = _io_result_T_1 ? _io_result_T_67 : _io_result_T_70; // @[FP16Add.scala 87:120]
  wire [15:0] _io_result_T_72 = _io_result_T_2 ? _io_result_T_63 : _io_result_T_71; // @[FP16Add.scala 87:25]
  wire [15:0] _GEN_3 = expA == expB ? _GEN_2 : _io_result_T_72; // @[FP16Add.scala 73:32 87:19]
  wire [15:0] _GEN_6 = expA > expB ? _io_result_T_18 : _GEN_3; // @[FP16Add.scala 69:24 72:19]
  wire [15:0] _GEN_7 = infFlagA | infFlagB ? _GEN_0 : _GEN_6; // @[FP16Add.scala 56:38]
  wire [15:0] _GEN_9 = zeroFlagA & ~zeroFlagB ? io_b : _GEN_7; // @[FP16Add.scala 53:41 55:17]
  wire [15:0] _GEN_11 = ~zeroFlagA & zeroFlagB ? io_a : _GEN_9; // @[FP16Add.scala 50:40 52:17]
  assign io_result = zeroFlagA & zeroFlagB ? 16'h0 : _GEN_11; // @[FP16Add.scala 46:32 48:17]
endmodule
