module FP16Add(
  input         clock,
  input         reset,
  input  [15:0] io_a,
  input  [15:0] io_b,
  output [15:0] io_result
);
  wire  signA = io_a[15]; // @[FP16Add.scala 13:18]
  wire [4:0] expA = io_a[14:10]; // @[FP16Add.scala 14:22]
  wire [9:0] sigA = io_a[9:0]; // @[FP16Add.scala 15:25]
  wire  signB = io_b[15]; // @[FP16Add.scala 13:18]
  wire [4:0] expB = io_b[14:10]; // @[FP16Add.scala 14:22]
  wire [9:0] sigB = io_b[9:0]; // @[FP16Add.scala 15:25]
  wire  _zeroFlagA_T = expA == 5'h0; // @[FP16Add.scala 38:24]
  wire  _zeroFlagA_T_1 = sigA == 10'h0; // @[FP16Add.scala 38:40]
  wire  zeroFlagA = expA == 5'h0 & sigA == 10'h0; // @[FP16Add.scala 38:32]
  wire  _zeroFlagB_T = expB == 5'h0; // @[FP16Add.scala 39:24]
  wire  _zeroFlagB_T_1 = sigB == 10'h0; // @[FP16Add.scala 39:40]
  wire  zeroFlagB = expB == 5'h0 & sigB == 10'h0; // @[FP16Add.scala 39:32]
  wire  infFlagA = expA == 5'h1f & _zeroFlagA_T_1; // @[FP16Add.scala 44:38]
  wire  infFlagB = expB == 5'h1f & _zeroFlagB_T_1; // @[FP16Add.scala 45:38]
  wire  subNormA = _zeroFlagA_T & sigA != 10'h0; // @[FP16Add.scala 47:31]
  wire  subNormB = _zeroFlagB_T & sigB != 10'h0; // @[FP16Add.scala 48:31]
  wire [15:0] _io_result_T = infFlagA ? io_a : io_b; // @[FP16Add.scala 72:25]
  wire [15:0] _GEN_0 = infFlagA & infFlagB & signA != signB ? 16'h7fff : _io_result_T; // @[FP16Add.scala 66:54 68:19 72:19]
  wire [9:0] _GEN_13 = {{5'd0}, expA}; // @[FP16Add.scala 74:49]
  wire [9:0] _GEN_14 = {{5'd0}, expB}; // @[FP16Add.scala 74:106]
  wire  _T_20 = ~signA; // @[FP16Add.scala 85:22]
  wire  _T_21 = ~signB; // @[FP16Add.scala 85:39]
  wire [10:0] _io_result_T_1 = {1'h1,sigA}; // @[Cat.scala 33:92]
  wire [10:0] _io_result_T_2 = {1'h1,sigB}; // @[Cat.scala 33:92]
  wire [11:0] _io_result_T_3 = _io_result_T_1 + _io_result_T_2; // @[FP16Add.scala 88:46]
  wire [4:0] _io_result_T_7 = expA + 5'h1; // @[FP16Add.scala 88:94]
  wire [15:0] _io_result_T_12 = {signA,_io_result_T_7,_io_result_T_3[10:1]}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_17 = {signA,expA,_io_result_T_3[9:0]}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_18 = _io_result_T_3[11] ? _io_result_T_12 : _io_result_T_17; // @[FP16Add.scala 88:29]
  wire  _io_result_T_19 = sigB >= sigA; // @[FP16Add.scala 91:35]
  wire [10:0] _io_result_T_23 = _io_result_T_2 - _io_result_T_1; // @[FP16Add.scala 91:75]
  wire [15:0] _io_result_T_25 = {1'h0,expB,_io_result_T_23[9:0]}; // @[Cat.scala 33:92]
  wire [10:0] _io_result_T_29 = _io_result_T_1 - _io_result_T_2; // @[FP16Add.scala 91:131]
  wire [15:0] _io_result_T_31 = {1'h1,expA,_io_result_T_29[9:0]}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_32 = sigB >= sigA ? _io_result_T_25 : _io_result_T_31; // @[FP16Add.scala 91:29]
  wire [15:0] _io_result_T_39 = {1'h1,expB,_io_result_T_23[9:0]}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_45 = {1'h0,expA,_io_result_T_29[9:0]}; // @[Cat.scala 33:92]
  wire [15:0] _io_result_T_46 = _io_result_T_19 ? _io_result_T_39 : _io_result_T_45; // @[FP16Add.scala 93:29]
  wire [15:0] _GEN_1 = _T_20 & signB ? _io_result_T_46 : _io_result_T_18; // @[FP16Add.scala 92:53 93:23 95:23]
  wire [15:0] _GEN_2 = signA & _T_21 ? _io_result_T_32 : _GEN_1; // @[FP16Add.scala 89:53 91:23]
  wire [15:0] _GEN_3 = ~signA & ~signB ? _io_result_T_18 : _GEN_2; // @[FP16Add.scala 85:47 88:23]
  wire [15:0] _GEN_5 = expA == expB ? _GEN_3 : 16'h0; // @[FP16Add.scala 82:29]
  wire [15:0] _GEN_7 = ~subNormA & ~subNormB ? _GEN_5 : 16'h0; // @[FP16Add.scala 79:34]
  wire [15:0] _GEN_8 = sigA == 10'h1f & _GEN_13 == 10'h3ff | sigB == 10'h1f & _GEN_14 == 10'h3ff ? 16'h7fff : _GEN_7; // @[FP16Add.scala 74:128 75:17]
  wire [15:0] _GEN_9 = infFlagA | infFlagB ? _GEN_0 : _GEN_8; // @[FP16Add.scala 64:38]
  wire [15:0] _GEN_10 = zeroFlagA & ~zeroFlagB ? io_b : _GEN_9; // @[FP16Add.scala 61:41 63:17]
  wire [15:0] _GEN_11 = ~zeroFlagA & zeroFlagB ? io_a : _GEN_10; // @[FP16Add.scala 58:40 60:17]
  assign io_result = zeroFlagA & zeroFlagB ? 16'h0 : _GEN_11; // @[FP16Add.scala 54:32 56:17]
endmodule
