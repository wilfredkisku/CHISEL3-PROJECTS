module INT8_MUL(
  input         clock,
  input         reset,
  input  [7:0]  io_inputA,
  input  [7:0]  io_inputB,
  output [15:0] io_output
);
  assign io_output = $signed(io_inputA) * $signed(io_inputB); // @[INT8_MUL.scala 12:26]
endmodule
