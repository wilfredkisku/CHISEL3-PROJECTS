module FP8_ADD(
  input        clock,
  input        reset,
  input  [7:0] io_inputA,
  input  [7:0] io_inputB,
  output [7:0] io_output
);
  wire  signA = io_inputA[7]; // @[FP8_ADD.scala 13:18]
  wire [4:0] expA = io_inputA[6:2]; // @[FP8_ADD.scala 14:22]
  wire [1:0] sigA = io_inputA[1:0]; // @[FP8_ADD.scala 15:25]
  wire  signB = io_inputB[7]; // @[FP8_ADD.scala 13:18]
  wire [4:0] expB = io_inputB[6:2]; // @[FP8_ADD.scala 14:22]
  wire [1:0] sigB = io_inputB[1:0]; // @[FP8_ADD.scala 15:25]
  wire  _infFlagA_T = expA == 5'h1f; // @[FP8_ADD.scala 24:23]
  wire  _infFlagA_T_1 = sigA == 2'h0; // @[FP8_ADD.scala 24:46]
  wire  infFlagA = expA == 5'h1f & sigA == 2'h0; // @[FP8_ADD.scala 24:38]
  wire  _infFlagB_T = expB == 5'h1f; // @[FP8_ADD.scala 25:23]
  wire  _infFlagB_T_1 = sigB == 2'h0; // @[FP8_ADD.scala 25:46]
  wire  infFlagB = expB == 5'h1f & sigB == 2'h0; // @[FP8_ADD.scala 25:38]
  wire  _zeroFlagA_T = expA == 5'h0; // @[FP8_ADD.scala 28:24]
  wire  zeroFlagA = expA == 5'h0 & _infFlagA_T_1; // @[FP8_ADD.scala 28:39]
  wire  _zeroFlagB_T = expB == 5'h0; // @[FP8_ADD.scala 29:24]
  wire  zeroFlagB = expB == 5'h0 & _infFlagB_T_1; // @[FP8_ADD.scala 29:39]
  wire  _nanFlagA_T_1 = sigA != 2'h0; // @[FP8_ADD.scala 32:46]
  wire  nanFlagA = _infFlagA_T & sigA != 2'h0; // @[FP8_ADD.scala 32:38]
  wire  _nanFlagB_T_1 = sigB != 2'h0; // @[FP8_ADD.scala 33:46]
  wire  nanFlagB = _infFlagB_T & sigB != 2'h0; // @[FP8_ADD.scala 33:38]
  wire  subFlagA = _zeroFlagA_T & _nanFlagA_T_1; // @[FP8_ADD.scala 36:38]
  wire  subFlagB = _zeroFlagB_T & _nanFlagB_T_1; // @[FP8_ADD.scala 37:38]
  wire [7:0] _io_output_T = zeroFlagA ? io_inputB : io_inputA; // @[FP8_ADD.scala 51:21]
  wire  _T_4 = signA != signB; // @[FP8_ADD.scala 54:42]
  wire [7:0] _io_output_T_1 = infFlagA ? io_inputA : io_inputB; // @[FP8_ADD.scala 57:23]
  wire [7:0] _GEN_0 = infFlagA & infFlagB & signA != signB ? 8'h7f : _io_output_T_1; // @[FP8_ADD.scala 54:53 55:17 57:17]
  wire [2:0] _ovrChk_a_T = {1'h1,sigA}; // @[Cat.scala 33:92]
  wire [2:0] _ovrChk_a_T_1 = {1'h1,sigB}; // @[Cat.scala 33:92]
  wire [4:0] _ovrChk_a_T_3 = expA - expB; // @[FP8_ADD.scala 82:64]
  wire [2:0] _ovrChk_a_T_4 = _ovrChk_a_T_1 >> _ovrChk_a_T_3; // @[FP8_ADD.scala 82:55]
  wire [3:0] _ovrChk_a_T_5 = _ovrChk_a_T + _ovrChk_a_T_4; // @[FP8_ADD.scala 82:36]
  wire [2:0] _ovrChk_s_T_6 = _ovrChk_a_T - _ovrChk_a_T_4; // @[FP8_ADD.scala 83:36]
  wire  _io_output_T_2 = ~signA; // @[FP8_ADD.scala 84:32]
  wire  _io_output_T_3 = ~signB; // @[FP8_ADD.scala 84:68]
  wire [4:0] _ovrChk_a_T_9 = expB - expA; // @[FP8_ADD.scala 87:64]
  wire [2:0] _ovrChk_a_T_10 = _ovrChk_a_T >> _ovrChk_a_T_9; // @[FP8_ADD.scala 87:55]
  wire [3:0] _ovrChk_a_T_11 = _ovrChk_a_T_1 + _ovrChk_a_T_10; // @[FP8_ADD.scala 87:36]
  wire [3:0] _GEN_3 = expB > expA ? _ovrChk_a_T_11 : _ovrChk_a_T_11; // @[FP8_ADD.scala 85:30 87:18 91:18]
  wire [3:0] _GEN_6 = expA > expB ? _ovrChk_a_T_5 : _GEN_3; // @[FP8_ADD.scala 80:24 82:18]
  wire [3:0] _GEN_9 = ~subFlagA & ~subFlagB ? _GEN_6 : 4'h0; // @[FP8_ADD.scala 43:12 71:39]
  wire [3:0] _GEN_13 = subFlagA & subFlagB ? 4'h0 : _GEN_9; // @[FP8_ADD.scala 43:12 63:31]
  wire [3:0] _GEN_16 = nanFlagA | nanFlagB ? 4'h0 : _GEN_13; // @[FP8_ADD.scala 43:12 59:35]
  wire [3:0] _GEN_19 = infFlagA | infFlagB ? 4'h0 : _GEN_16; // @[FP8_ADD.scala 43:12 52:35]
  wire [3:0] _GEN_22 = zeroFlagA | zeroFlagB ? 4'h0 : _GEN_19; // @[FP8_ADD.scala 43:12 50:37]
  wire [3:0] ovrChk_a = zeroFlagA & zeroFlagB ? 4'h0 : _GEN_22; // @[FP8_ADD.scala 43:12 47:32]
  wire [2:0] _ovrChk_s_T_13 = _ovrChk_a_T_1 - _ovrChk_a_T_10; // @[FP8_ADD.scala 88:36]
  wire [2:0] _GEN_4 = expB > expA ? _ovrChk_s_T_13 : _ovrChk_s_T_13; // @[FP8_ADD.scala 85:30 88:18 92:18]
  wire [2:0] _GEN_7 = expA > expB ? _ovrChk_s_T_6 : _GEN_4; // @[FP8_ADD.scala 80:24 83:18]
  wire [2:0] _GEN_10 = ~subFlagA & ~subFlagB ? _GEN_7 : 3'h0; // @[FP8_ADD.scala 44:12 71:39]
  wire [2:0] _GEN_14 = subFlagA & subFlagB ? 3'h0 : _GEN_10; // @[FP8_ADD.scala 44:12 63:31]
  wire [2:0] _GEN_17 = nanFlagA | nanFlagB ? 3'h0 : _GEN_14; // @[FP8_ADD.scala 44:12 59:35]
  wire [2:0] _GEN_20 = infFlagA | infFlagB ? 3'h0 : _GEN_17; // @[FP8_ADD.scala 44:12 52:35]
  wire [2:0] _GEN_23 = zeroFlagA | zeroFlagB ? 3'h0 : _GEN_20; // @[FP8_ADD.scala 44:12 50:37]
  wire [2:0] _GEN_26 = zeroFlagA & zeroFlagB ? 3'h0 : _GEN_23; // @[FP8_ADD.scala 44:12 47:32]
  wire [3:0] ovrChk_s = {{1'd0}, _GEN_26}; // @[FP8_ADD.scala 41:22]
  wire [1:0] _io_output_T_6 = ~signB ? ovrChk_a[1:0] : ovrChk_s[1:0]; // @[FP8_ADD.scala 84:61]
  wire [7:0] _io_output_T_7 = {signA,expA,_io_output_T_6}; // @[Cat.scala 33:92]
  wire [1:0] _io_output_T_11 = ~signB ? ovrChk_s[1:0] : ovrChk_a[1:0]; // @[FP8_ADD.scala 84:129]
  wire [7:0] _io_output_T_12 = {signA,expA,_io_output_T_11}; // @[Cat.scala 33:92]
  wire [7:0] _io_output_T_13 = ~signA ? _io_output_T_7 : _io_output_T_12; // @[FP8_ADD.scala 84:25]
  wire [1:0] _io_output_T_18 = _io_output_T_2 ? ovrChk_s[1:0] : ovrChk_a[1:0]; // @[FP8_ADD.scala 89:61]
  wire [7:0] _io_output_T_19 = {signB,expB,_io_output_T_18}; // @[Cat.scala 33:92]
  wire [1:0] _io_output_T_23 = _io_output_T_2 ? ovrChk_a[1:0] : ovrChk_s[1:0]; // @[FP8_ADD.scala 89:129]
  wire [7:0] _io_output_T_24 = {signB,expB,_io_output_T_23}; // @[Cat.scala 33:92]
  wire [7:0] _io_output_T_25 = _io_output_T_3 ? _io_output_T_19 : _io_output_T_24; // @[FP8_ADD.scala 89:25]
  wire [4:0] _GEN_27 = {{4'd0}, ovrChk_a[3]}; // @[FP8_ADD.scala 99:66]
  wire [4:0] _io_output_T_29 = expA + _GEN_27; // @[FP8_ADD.scala 99:66]
  wire [3:0] _io_output_T_31 = ovrChk_a >> ovrChk_a[3]; // @[FP8_ADD.scala 99:91]
  wire [7:0] _io_output_T_33 = {signA,_io_output_T_29,_io_output_T_31[1:0]}; // @[Cat.scala 33:92]
  wire [7:0] _io_output_T_34 = _T_4 ? 8'h0 : _io_output_T_33; // @[FP8_ADD.scala 99:27]
  wire [7:0] _GEN_1 = sigB > sigA ? 8'h0 : _io_output_T_34; // @[FP8_ADD.scala 96:32 97:21 99:21]
  wire [7:0] _GEN_2 = sigA > sigB ? 8'h0 : _GEN_1; // @[FP8_ADD.scala 94:26 95:21]
  wire [7:0] _GEN_5 = expB > expA ? _io_output_T_25 : _GEN_2; // @[FP8_ADD.scala 85:30 89:19]
  wire [7:0] _GEN_8 = expA > expB ? _io_output_T_13 : _GEN_5; // @[FP8_ADD.scala 80:24 84:19]
  wire [7:0] _GEN_11 = ~subFlagA & ~subFlagB ? _GEN_8 : 8'h0; // @[FP8_ADD.scala 109:17 71:39]
  wire [7:0] _GEN_12 = subFlagA & subFlagB ? 8'h0 : _GEN_11; // @[FP8_ADD.scala 63:31 67:17]
  wire [7:0] _GEN_15 = nanFlagA | nanFlagB ? 8'h7f : _GEN_12; // @[FP8_ADD.scala 59:35 60:15]
  wire [7:0] _GEN_18 = infFlagA | infFlagB ? _GEN_0 : _GEN_15; // @[FP8_ADD.scala 52:35]
  wire [7:0] _GEN_21 = zeroFlagA | zeroFlagB ? _io_output_T : _GEN_18; // @[FP8_ADD.scala 50:37 51:15]
  assign io_output = zeroFlagA & zeroFlagB ? 8'h0 : _GEN_21; // @[FP8_ADD.scala 47:32 49:15]
endmodule
