module BufferAMSNew(
  input        clock,
  input        reset,
  input  [7:0] io_adcValues_0,
  input  [7:0] io_adcValues_1,
  input  [7:0] io_adcValues_2,
  input  [7:0] io_adcValues_3,
  input  [7:0] io_adcValues_4,
  input  [7:0] io_adcValues_5,
  input  [7:0] io_adcValues_6,
  input  [7:0] io_adcValues_7,
  input  [7:0] io_adcValues_8,
  input  [7:0] io_adcValues_9,
  input  [7:0] io_adcValues_10,
  input  [7:0] io_adcValues_11,
  input  [7:0] io_adcValues_12,
  input  [7:0] io_adcValues_13,
  input  [7:0] io_adcValues_14,
  input  [7:0] io_adcValues_15,
  input  [7:0] io_adcValues_16,
  input  [7:0] io_adcValues_17,
  input  [7:0] io_adcValues_18,
  input  [7:0] io_adcValues_19,
  input  [7:0] io_adcValues_20,
  input  [7:0] io_adcValues_21,
  input  [7:0] io_adcValues_22,
  input  [7:0] io_adcValues_23,
  input  [7:0] io_adcValues_24,
  input  [7:0] io_adcValues_25,
  input  [7:0] io_adcValues_26,
  input  [7:0] io_adcValues_27,
  input  [7:0] io_adcValues_28,
  input  [7:0] io_adcValues_29,
  input  [7:0] io_adcValues_30,
  input  [7:0] io_adcValues_31,
  input  [7:0] io_adcValues_32,
  input  [7:0] io_adcValues_33,
  input  [7:0] io_adcValues_34,
  input  [7:0] io_adcValues_35,
  input  [7:0] io_adcValues_36,
  input  [7:0] io_adcValues_37,
  input  [7:0] io_adcValues_38,
  input  [7:0] io_adcValues_39,
  input  [7:0] io_adcValues_40,
  input  [7:0] io_adcValues_41,
  input  [7:0] io_adcValues_42,
  input  [7:0] io_adcValues_43,
  input  [7:0] io_adcValues_44,
  input  [7:0] io_adcValues_45,
  input  [7:0] io_adcValues_46,
  input  [7:0] io_adcValues_47,
  input  [7:0] io_adcValues_48,
  input  [7:0] io_adcValues_49,
  input  [7:0] io_adcValues_50,
  input  [7:0] io_adcValues_51,
  input  [7:0] io_adcValues_52,
  input  [7:0] io_adcValues_53,
  input  [7:0] io_adcValues_54,
  input  [7:0] io_adcValues_55,
  input  [7:0] io_adcValues_56,
  input  [7:0] io_adcValues_57,
  input  [7:0] io_adcValues_58,
  input  [7:0] io_adcValues_59,
  input  [7:0] io_adcValues_60,
  input  [7:0] io_adcValues_61,
  input  [7:0] io_adcValues_62,
  input  [7:0] io_adcValues_63,
  input  [7:0] io_adcValues_64,
  input  [7:0] io_adcValues_65,
  input  [7:0] io_adcValues_66,
  input  [7:0] io_adcValues_67,
  input  [7:0] io_adcValues_68,
  input  [7:0] io_adcValues_69,
  input  [7:0] io_adcValues_70,
  input  [7:0] io_adcValues_71,
  input  [7:0] io_adcValues_72,
  input  [7:0] io_adcValues_73,
  input  [7:0] io_adcValues_74,
  input  [7:0] io_adcValues_75,
  input  [7:0] io_adcValues_76,
  input  [7:0] io_adcValues_77,
  input  [7:0] io_adcValues_78,
  input  [7:0] io_adcValues_79,
  input  [7:0] io_adcValues_80,
  input  [7:0] io_adcValues_81,
  input  [7:0] io_adcValues_82,
  input  [7:0] io_adcValues_83,
  input  [7:0] io_adcValues_84,
  input  [7:0] io_adcValues_85,
  input  [7:0] io_adcValues_86,
  input  [7:0] io_adcValues_87,
  input  [7:0] io_adcValues_88,
  input  [7:0] io_adcValues_89,
  input  [7:0] io_adcValues_90,
  input  [7:0] io_adcValues_91,
  input  [7:0] io_adcValues_92,
  input  [7:0] io_adcValues_93,
  input  [7:0] io_adcValues_94,
  input  [7:0] io_adcValues_95,
  input  [7:0] io_adcValues_96,
  input  [7:0] io_adcValues_97,
  input  [7:0] io_adcValues_98,
  input  [7:0] io_adcValues_99,
  input  [7:0] io_adcValues_100,
  input  [7:0] io_adcValues_101,
  input  [7:0] io_adcValues_102,
  input  [7:0] io_adcValues_103,
  input  [7:0] io_adcValues_104,
  input  [7:0] io_adcValues_105,
  input  [7:0] io_adcValues_106,
  input  [7:0] io_adcValues_107,
  input  [7:0] io_adcValues_108,
  input  [7:0] io_adcValues_109,
  input  [7:0] io_adcValues_110,
  input  [7:0] io_adcValues_111,
  input  [7:0] io_adcValues_112,
  input  [7:0] io_adcValues_113,
  input  [7:0] io_adcValues_114,
  input  [7:0] io_adcValues_115,
  input  [7:0] io_adcValues_116,
  input  [7:0] io_adcValues_117,
  input  [7:0] io_adcValues_118,
  input  [7:0] io_adcValues_119,
  input  [7:0] io_adcValues_120,
  input  [7:0] io_adcValues_121,
  input  [7:0] io_adcValues_122,
  input  [7:0] io_adcValues_123,
  input  [7:0] io_adcValues_124,
  input  [7:0] io_adcValues_125,
  input  [7:0] io_adcValues_126,
  input  [7:0] io_adcValues_127,
  output [7:0] io_zeroSums_0,
  output [7:0] io_zeroSums_1,
  output [7:0] io_zeroSums_2,
  output [7:0] io_zeroSums_3,
  output [7:0] io_zeroSums_4,
  output [7:0] io_zeroSums_5,
  output [7:0] io_zeroSums_6,
  output [7:0] io_zeroSums_7,
  output [3:0] io_indicesOut_0,
  output [3:0] io_indicesOut_1,
  output [3:0] io_indicesOut_2,
  output [3:0] io_indicesOut_3,
  output [3:0] io_indicesOut_4,
  output [3:0] io_indicesOut_5,
  output [3:0] io_indicesOut_6,
  output [3:0] io_indicesOut_7,
  output [7:0] io_frameOut_0,
  output [7:0] io_frameOut_1,
  output [7:0] io_frameOut_2,
  output [7:0] io_frameOut_3,
  output [7:0] io_frameOut_4,
  output [7:0] io_frameOut_5,
  output [7:0] io_frameOut_6,
  output [7:0] io_frameOut_7,
  output [7:0] io_frameOut_8,
  output [7:0] io_frameOut_9,
  output [7:0] io_frameOut_10,
  output [7:0] io_frameOut_11,
  output [7:0] io_frameOut_12,
  output [7:0] io_frameOut_13,
  output [7:0] io_frameOut_14,
  output [7:0] io_frameOut_15,
  output [7:0] io_frameOut_16,
  output [7:0] io_frameOut_17,
  output [7:0] io_frameOut_18,
  output [7:0] io_frameOut_19,
  output [7:0] io_frameOut_20,
  output [7:0] io_frameOut_21,
  output [7:0] io_frameOut_22,
  output [7:0] io_frameOut_23,
  output [7:0] io_frameOut_24,
  output [7:0] io_frameOut_25,
  output [7:0] io_frameOut_26,
  output [7:0] io_frameOut_27,
  output [7:0] io_frameOut_28,
  output [7:0] io_frameOut_29,
  output [7:0] io_frameOut_30,
  output [7:0] io_frameOut_31,
  output [7:0] io_frameOut_32,
  output [7:0] io_frameOut_33,
  output [7:0] io_frameOut_34,
  output [7:0] io_frameOut_35,
  output [7:0] io_frameOut_36,
  output [7:0] io_frameOut_37,
  output [7:0] io_frameOut_38,
  output [7:0] io_frameOut_39,
  output [7:0] io_frameOut_40,
  output [7:0] io_frameOut_41,
  output [7:0] io_frameOut_42,
  output [7:0] io_frameOut_43,
  output [7:0] io_frameOut_44,
  output [7:0] io_frameOut_45,
  output [7:0] io_frameOut_46,
  output [7:0] io_frameOut_47,
  output [7:0] io_frameOut_48,
  output [7:0] io_frameOut_49,
  output [7:0] io_frameOut_50,
  output [7:0] io_frameOut_51,
  output [7:0] io_frameOut_52,
  output [7:0] io_frameOut_53,
  output [7:0] io_frameOut_54,
  output [7:0] io_frameOut_55,
  output [7:0] io_frameOut_56,
  output [7:0] io_frameOut_57,
  output [7:0] io_frameOut_58,
  output [7:0] io_frameOut_59,
  output [7:0] io_frameOut_60,
  output [7:0] io_frameOut_61,
  output [7:0] io_frameOut_62,
  output [7:0] io_frameOut_63,
  output [7:0] io_frameOut_64,
  output [7:0] io_frameOut_65,
  output [7:0] io_frameOut_66,
  output [7:0] io_frameOut_67,
  output [7:0] io_frameOut_68,
  output [7:0] io_frameOut_69,
  output [7:0] io_frameOut_70,
  output [7:0] io_frameOut_71,
  output [7:0] io_frameOut_72,
  output [7:0] io_frameOut_73,
  output [7:0] io_frameOut_74,
  output [7:0] io_frameOut_75,
  output [7:0] io_frameOut_76,
  output [7:0] io_frameOut_77,
  output [7:0] io_frameOut_78,
  output [7:0] io_frameOut_79,
  output [7:0] io_frameOut_80,
  output [7:0] io_frameOut_81,
  output [7:0] io_frameOut_82,
  output [7:0] io_frameOut_83,
  output [7:0] io_frameOut_84,
  output [7:0] io_frameOut_85,
  output [7:0] io_frameOut_86,
  output [7:0] io_frameOut_87,
  output [7:0] io_frameOut_88,
  output [7:0] io_frameOut_89,
  output [7:0] io_frameOut_90,
  output [7:0] io_frameOut_91,
  output [7:0] io_frameOut_92,
  output [7:0] io_frameOut_93,
  output [7:0] io_frameOut_94,
  output [7:0] io_frameOut_95,
  output [7:0] io_frameOut_96,
  output [7:0] io_frameOut_97,
  output [7:0] io_frameOut_98,
  output [7:0] io_frameOut_99,
  output [7:0] io_frameOut_100,
  output [7:0] io_frameOut_101,
  output [7:0] io_frameOut_102,
  output [7:0] io_frameOut_103,
  output [7:0] io_frameOut_104,
  output [7:0] io_frameOut_105,
  output [7:0] io_frameOut_106,
  output [7:0] io_frameOut_107,
  output [7:0] io_frameOut_108,
  output [7:0] io_frameOut_109,
  output [7:0] io_frameOut_110,
  output [7:0] io_frameOut_111,
  output [7:0] io_frameOut_112,
  output [7:0] io_frameOut_113,
  output [7:0] io_frameOut_114,
  output [7:0] io_frameOut_115,
  output [7:0] io_frameOut_116,
  output [7:0] io_frameOut_117,
  output [7:0] io_frameOut_118,
  output [7:0] io_frameOut_119,
  output [7:0] io_frameOut_120,
  output [7:0] io_frameOut_121,
  output [7:0] io_frameOut_122,
  output [7:0] io_frameOut_123,
  output [7:0] io_frameOut_124,
  output [7:0] io_frameOut_125,
  output [7:0] io_frameOut_126,
  output [7:0] io_frameOut_127
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
  reg [31:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1560;
  reg [31:0] _RAND_1561;
  reg [31:0] _RAND_1562;
  reg [31:0] _RAND_1563;
  reg [31:0] _RAND_1564;
  reg [31:0] _RAND_1565;
  reg [31:0] _RAND_1566;
  reg [31:0] _RAND_1567;
  reg [31:0] _RAND_1568;
  reg [31:0] _RAND_1569;
  reg [31:0] _RAND_1570;
  reg [31:0] _RAND_1571;
  reg [31:0] _RAND_1572;
  reg [31:0] _RAND_1573;
  reg [31:0] _RAND_1574;
  reg [31:0] _RAND_1575;
  reg [31:0] _RAND_1576;
  reg [31:0] _RAND_1577;
  reg [31:0] _RAND_1578;
  reg [31:0] _RAND_1579;
  reg [31:0] _RAND_1580;
  reg [31:0] _RAND_1581;
  reg [31:0] _RAND_1582;
  reg [31:0] _RAND_1583;
  reg [31:0] _RAND_1584;
  reg [31:0] _RAND_1585;
  reg [31:0] _RAND_1586;
  reg [31:0] _RAND_1587;
  reg [31:0] _RAND_1588;
  reg [31:0] _RAND_1589;
  reg [31:0] _RAND_1590;
  reg [31:0] _RAND_1591;
  reg [31:0] _RAND_1592;
  reg [31:0] _RAND_1593;
  reg [31:0] _RAND_1594;
  reg [31:0] _RAND_1595;
  reg [31:0] _RAND_1596;
  reg [31:0] _RAND_1597;
  reg [31:0] _RAND_1598;
  reg [31:0] _RAND_1599;
  reg [31:0] _RAND_1600;
  reg [31:0] _RAND_1601;
  reg [31:0] _RAND_1602;
  reg [31:0] _RAND_1603;
  reg [31:0] _RAND_1604;
  reg [31:0] _RAND_1605;
  reg [31:0] _RAND_1606;
  reg [31:0] _RAND_1607;
  reg [31:0] _RAND_1608;
  reg [31:0] _RAND_1609;
  reg [31:0] _RAND_1610;
  reg [31:0] _RAND_1611;
  reg [31:0] _RAND_1612;
  reg [31:0] _RAND_1613;
  reg [31:0] _RAND_1614;
  reg [31:0] _RAND_1615;
  reg [31:0] _RAND_1616;
  reg [31:0] _RAND_1617;
  reg [31:0] _RAND_1618;
  reg [31:0] _RAND_1619;
  reg [31:0] _RAND_1620;
  reg [31:0] _RAND_1621;
  reg [31:0] _RAND_1622;
  reg [31:0] _RAND_1623;
  reg [31:0] _RAND_1624;
  reg [31:0] _RAND_1625;
  reg [31:0] _RAND_1626;
  reg [31:0] _RAND_1627;
  reg [31:0] _RAND_1628;
  reg [31:0] _RAND_1629;
  reg [31:0] _RAND_1630;
  reg [31:0] _RAND_1631;
  reg [31:0] _RAND_1632;
  reg [31:0] _RAND_1633;
  reg [31:0] _RAND_1634;
  reg [31:0] _RAND_1635;
  reg [31:0] _RAND_1636;
  reg [31:0] _RAND_1637;
  reg [31:0] _RAND_1638;
  reg [31:0] _RAND_1639;
  reg [31:0] _RAND_1640;
  reg [31:0] _RAND_1641;
  reg [31:0] _RAND_1642;
  reg [31:0] _RAND_1643;
  reg [31:0] _RAND_1644;
  reg [31:0] _RAND_1645;
  reg [31:0] _RAND_1646;
  reg [31:0] _RAND_1647;
  reg [31:0] _RAND_1648;
  reg [31:0] _RAND_1649;
  reg [31:0] _RAND_1650;
  reg [31:0] _RAND_1651;
  reg [31:0] _RAND_1652;
  reg [31:0] _RAND_1653;
  reg [31:0] _RAND_1654;
  reg [31:0] _RAND_1655;
  reg [31:0] _RAND_1656;
  reg [31:0] _RAND_1657;
  reg [31:0] _RAND_1658;
  reg [31:0] _RAND_1659;
  reg [31:0] _RAND_1660;
  reg [31:0] _RAND_1661;
  reg [31:0] _RAND_1662;
  reg [31:0] _RAND_1663;
  reg [31:0] _RAND_1664;
  reg [31:0] _RAND_1665;
  reg [31:0] _RAND_1666;
  reg [31:0] _RAND_1667;
  reg [31:0] _RAND_1668;
  reg [31:0] _RAND_1669;
  reg [31:0] _RAND_1670;
  reg [31:0] _RAND_1671;
  reg [31:0] _RAND_1672;
  reg [31:0] _RAND_1673;
  reg [31:0] _RAND_1674;
  reg [31:0] _RAND_1675;
  reg [31:0] _RAND_1676;
  reg [31:0] _RAND_1677;
  reg [31:0] _RAND_1678;
  reg [31:0] _RAND_1679;
  reg [31:0] _RAND_1680;
  reg [31:0] _RAND_1681;
  reg [31:0] _RAND_1682;
  reg [31:0] _RAND_1683;
  reg [31:0] _RAND_1684;
  reg [31:0] _RAND_1685;
  reg [31:0] _RAND_1686;
  reg [31:0] _RAND_1687;
  reg [31:0] _RAND_1688;
  reg [31:0] _RAND_1689;
  reg [31:0] _RAND_1690;
  reg [31:0] _RAND_1691;
  reg [31:0] _RAND_1692;
  reg [31:0] _RAND_1693;
  reg [31:0] _RAND_1694;
  reg [31:0] _RAND_1695;
  reg [31:0] _RAND_1696;
  reg [31:0] _RAND_1697;
  reg [31:0] _RAND_1698;
  reg [31:0] _RAND_1699;
  reg [31:0] _RAND_1700;
  reg [31:0] _RAND_1701;
  reg [31:0] _RAND_1702;
  reg [31:0] _RAND_1703;
  reg [31:0] _RAND_1704;
  reg [31:0] _RAND_1705;
  reg [31:0] _RAND_1706;
  reg [31:0] _RAND_1707;
  reg [31:0] _RAND_1708;
  reg [31:0] _RAND_1709;
  reg [31:0] _RAND_1710;
  reg [31:0] _RAND_1711;
  reg [31:0] _RAND_1712;
  reg [31:0] _RAND_1713;
  reg [31:0] _RAND_1714;
  reg [31:0] _RAND_1715;
  reg [31:0] _RAND_1716;
  reg [31:0] _RAND_1717;
  reg [31:0] _RAND_1718;
  reg [31:0] _RAND_1719;
  reg [31:0] _RAND_1720;
  reg [31:0] _RAND_1721;
  reg [31:0] _RAND_1722;
  reg [31:0] _RAND_1723;
  reg [31:0] _RAND_1724;
  reg [31:0] _RAND_1725;
  reg [31:0] _RAND_1726;
  reg [31:0] _RAND_1727;
  reg [31:0] _RAND_1728;
  reg [31:0] _RAND_1729;
  reg [31:0] _RAND_1730;
  reg [31:0] _RAND_1731;
  reg [31:0] _RAND_1732;
  reg [31:0] _RAND_1733;
  reg [31:0] _RAND_1734;
  reg [31:0] _RAND_1735;
  reg [31:0] _RAND_1736;
  reg [31:0] _RAND_1737;
  reg [31:0] _RAND_1738;
  reg [31:0] _RAND_1739;
  reg [31:0] _RAND_1740;
  reg [31:0] _RAND_1741;
  reg [31:0] _RAND_1742;
  reg [31:0] _RAND_1743;
  reg [31:0] _RAND_1744;
  reg [31:0] _RAND_1745;
  reg [31:0] _RAND_1746;
  reg [31:0] _RAND_1747;
  reg [31:0] _RAND_1748;
  reg [31:0] _RAND_1749;
  reg [31:0] _RAND_1750;
  reg [31:0] _RAND_1751;
  reg [31:0] _RAND_1752;
  reg [31:0] _RAND_1753;
  reg [31:0] _RAND_1754;
  reg [31:0] _RAND_1755;
  reg [31:0] _RAND_1756;
  reg [31:0] _RAND_1757;
  reg [31:0] _RAND_1758;
  reg [31:0] _RAND_1759;
  reg [31:0] _RAND_1760;
  reg [31:0] _RAND_1761;
  reg [31:0] _RAND_1762;
  reg [31:0] _RAND_1763;
  reg [31:0] _RAND_1764;
  reg [31:0] _RAND_1765;
  reg [31:0] _RAND_1766;
  reg [31:0] _RAND_1767;
  reg [31:0] _RAND_1768;
  reg [31:0] _RAND_1769;
  reg [31:0] _RAND_1770;
  reg [31:0] _RAND_1771;
  reg [31:0] _RAND_1772;
  reg [31:0] _RAND_1773;
  reg [31:0] _RAND_1774;
  reg [31:0] _RAND_1775;
  reg [31:0] _RAND_1776;
  reg [31:0] _RAND_1777;
  reg [31:0] _RAND_1778;
  reg [31:0] _RAND_1779;
  reg [31:0] _RAND_1780;
  reg [31:0] _RAND_1781;
  reg [31:0] _RAND_1782;
  reg [31:0] _RAND_1783;
  reg [31:0] _RAND_1784;
  reg [31:0] _RAND_1785;
  reg [31:0] _RAND_1786;
  reg [31:0] _RAND_1787;
  reg [31:0] _RAND_1788;
  reg [31:0] _RAND_1789;
  reg [31:0] _RAND_1790;
  reg [31:0] _RAND_1791;
  reg [31:0] _RAND_1792;
  reg [31:0] _RAND_1793;
  reg [31:0] _RAND_1794;
  reg [31:0] _RAND_1795;
  reg [31:0] _RAND_1796;
  reg [31:0] _RAND_1797;
  reg [31:0] _RAND_1798;
  reg [31:0] _RAND_1799;
  reg [31:0] _RAND_1800;
  reg [31:0] _RAND_1801;
  reg [31:0] _RAND_1802;
  reg [31:0] _RAND_1803;
  reg [31:0] _RAND_1804;
  reg [31:0] _RAND_1805;
  reg [31:0] _RAND_1806;
  reg [31:0] _RAND_1807;
  reg [31:0] _RAND_1808;
  reg [31:0] _RAND_1809;
  reg [31:0] _RAND_1810;
  reg [31:0] _RAND_1811;
  reg [31:0] _RAND_1812;
  reg [31:0] _RAND_1813;
  reg [31:0] _RAND_1814;
  reg [31:0] _RAND_1815;
  reg [31:0] _RAND_1816;
  reg [31:0] _RAND_1817;
  reg [31:0] _RAND_1818;
  reg [31:0] _RAND_1819;
  reg [31:0] _RAND_1820;
  reg [31:0] _RAND_1821;
  reg [31:0] _RAND_1822;
  reg [31:0] _RAND_1823;
  reg [31:0] _RAND_1824;
  reg [31:0] _RAND_1825;
  reg [31:0] _RAND_1826;
  reg [31:0] _RAND_1827;
  reg [31:0] _RAND_1828;
  reg [31:0] _RAND_1829;
  reg [31:0] _RAND_1830;
  reg [31:0] _RAND_1831;
  reg [31:0] _RAND_1832;
  reg [31:0] _RAND_1833;
  reg [31:0] _RAND_1834;
  reg [31:0] _RAND_1835;
  reg [31:0] _RAND_1836;
  reg [31:0] _RAND_1837;
  reg [31:0] _RAND_1838;
  reg [31:0] _RAND_1839;
  reg [31:0] _RAND_1840;
  reg [31:0] _RAND_1841;
  reg [31:0] _RAND_1842;
  reg [31:0] _RAND_1843;
  reg [31:0] _RAND_1844;
  reg [31:0] _RAND_1845;
  reg [31:0] _RAND_1846;
  reg [31:0] _RAND_1847;
  reg [31:0] _RAND_1848;
  reg [31:0] _RAND_1849;
  reg [31:0] _RAND_1850;
  reg [31:0] _RAND_1851;
  reg [31:0] _RAND_1852;
  reg [31:0] _RAND_1853;
  reg [31:0] _RAND_1854;
  reg [31:0] _RAND_1855;
  reg [31:0] _RAND_1856;
  reg [31:0] _RAND_1857;
  reg [31:0] _RAND_1858;
  reg [31:0] _RAND_1859;
  reg [31:0] _RAND_1860;
  reg [31:0] _RAND_1861;
  reg [31:0] _RAND_1862;
  reg [31:0] _RAND_1863;
  reg [31:0] _RAND_1864;
  reg [31:0] _RAND_1865;
  reg [31:0] _RAND_1866;
  reg [31:0] _RAND_1867;
  reg [31:0] _RAND_1868;
  reg [31:0] _RAND_1869;
  reg [31:0] _RAND_1870;
  reg [31:0] _RAND_1871;
  reg [31:0] _RAND_1872;
  reg [31:0] _RAND_1873;
  reg [31:0] _RAND_1874;
  reg [31:0] _RAND_1875;
  reg [31:0] _RAND_1876;
  reg [31:0] _RAND_1877;
  reg [31:0] _RAND_1878;
  reg [31:0] _RAND_1879;
  reg [31:0] _RAND_1880;
  reg [31:0] _RAND_1881;
  reg [31:0] _RAND_1882;
  reg [31:0] _RAND_1883;
  reg [31:0] _RAND_1884;
  reg [31:0] _RAND_1885;
  reg [31:0] _RAND_1886;
  reg [31:0] _RAND_1887;
  reg [31:0] _RAND_1888;
  reg [31:0] _RAND_1889;
  reg [31:0] _RAND_1890;
  reg [31:0] _RAND_1891;
  reg [31:0] _RAND_1892;
  reg [31:0] _RAND_1893;
  reg [31:0] _RAND_1894;
  reg [31:0] _RAND_1895;
  reg [31:0] _RAND_1896;
  reg [31:0] _RAND_1897;
  reg [31:0] _RAND_1898;
  reg [31:0] _RAND_1899;
  reg [31:0] _RAND_1900;
  reg [31:0] _RAND_1901;
  reg [31:0] _RAND_1902;
  reg [31:0] _RAND_1903;
  reg [31:0] _RAND_1904;
  reg [31:0] _RAND_1905;
  reg [31:0] _RAND_1906;
  reg [31:0] _RAND_1907;
  reg [31:0] _RAND_1908;
  reg [31:0] _RAND_1909;
  reg [31:0] _RAND_1910;
  reg [31:0] _RAND_1911;
  reg [31:0] _RAND_1912;
  reg [31:0] _RAND_1913;
  reg [31:0] _RAND_1914;
  reg [31:0] _RAND_1915;
  reg [31:0] _RAND_1916;
  reg [31:0] _RAND_1917;
  reg [31:0] _RAND_1918;
  reg [31:0] _RAND_1919;
  reg [31:0] _RAND_1920;
  reg [31:0] _RAND_1921;
  reg [31:0] _RAND_1922;
  reg [31:0] _RAND_1923;
  reg [31:0] _RAND_1924;
  reg [31:0] _RAND_1925;
  reg [31:0] _RAND_1926;
  reg [31:0] _RAND_1927;
  reg [31:0] _RAND_1928;
  reg [31:0] _RAND_1929;
  reg [31:0] _RAND_1930;
  reg [31:0] _RAND_1931;
  reg [31:0] _RAND_1932;
  reg [31:0] _RAND_1933;
  reg [31:0] _RAND_1934;
  reg [31:0] _RAND_1935;
  reg [31:0] _RAND_1936;
  reg [31:0] _RAND_1937;
  reg [31:0] _RAND_1938;
  reg [31:0] _RAND_1939;
  reg [31:0] _RAND_1940;
  reg [31:0] _RAND_1941;
  reg [31:0] _RAND_1942;
  reg [31:0] _RAND_1943;
  reg [31:0] _RAND_1944;
  reg [31:0] _RAND_1945;
  reg [31:0] _RAND_1946;
  reg [31:0] _RAND_1947;
  reg [31:0] _RAND_1948;
  reg [31:0] _RAND_1949;
  reg [31:0] _RAND_1950;
  reg [31:0] _RAND_1951;
  reg [31:0] _RAND_1952;
  reg [31:0] _RAND_1953;
  reg [31:0] _RAND_1954;
  reg [31:0] _RAND_1955;
  reg [31:0] _RAND_1956;
  reg [31:0] _RAND_1957;
  reg [31:0] _RAND_1958;
  reg [31:0] _RAND_1959;
  reg [31:0] _RAND_1960;
  reg [31:0] _RAND_1961;
  reg [31:0] _RAND_1962;
  reg [31:0] _RAND_1963;
  reg [31:0] _RAND_1964;
  reg [31:0] _RAND_1965;
  reg [31:0] _RAND_1966;
  reg [31:0] _RAND_1967;
  reg [31:0] _RAND_1968;
  reg [31:0] _RAND_1969;
  reg [31:0] _RAND_1970;
  reg [31:0] _RAND_1971;
  reg [31:0] _RAND_1972;
  reg [31:0] _RAND_1973;
  reg [31:0] _RAND_1974;
  reg [31:0] _RAND_1975;
  reg [31:0] _RAND_1976;
  reg [31:0] _RAND_1977;
  reg [31:0] _RAND_1978;
  reg [31:0] _RAND_1979;
  reg [31:0] _RAND_1980;
  reg [31:0] _RAND_1981;
  reg [31:0] _RAND_1982;
  reg [31:0] _RAND_1983;
  reg [31:0] _RAND_1984;
  reg [31:0] _RAND_1985;
  reg [31:0] _RAND_1986;
  reg [31:0] _RAND_1987;
  reg [31:0] _RAND_1988;
  reg [31:0] _RAND_1989;
  reg [31:0] _RAND_1990;
  reg [31:0] _RAND_1991;
  reg [31:0] _RAND_1992;
  reg [31:0] _RAND_1993;
  reg [31:0] _RAND_1994;
  reg [31:0] _RAND_1995;
  reg [31:0] _RAND_1996;
  reg [31:0] _RAND_1997;
  reg [31:0] _RAND_1998;
  reg [31:0] _RAND_1999;
  reg [31:0] _RAND_2000;
  reg [31:0] _RAND_2001;
  reg [31:0] _RAND_2002;
  reg [31:0] _RAND_2003;
  reg [31:0] _RAND_2004;
  reg [31:0] _RAND_2005;
  reg [31:0] _RAND_2006;
  reg [31:0] _RAND_2007;
  reg [31:0] _RAND_2008;
  reg [31:0] _RAND_2009;
  reg [31:0] _RAND_2010;
  reg [31:0] _RAND_2011;
  reg [31:0] _RAND_2012;
  reg [31:0] _RAND_2013;
  reg [31:0] _RAND_2014;
  reg [31:0] _RAND_2015;
  reg [31:0] _RAND_2016;
  reg [31:0] _RAND_2017;
  reg [31:0] _RAND_2018;
  reg [31:0] _RAND_2019;
  reg [31:0] _RAND_2020;
  reg [31:0] _RAND_2021;
  reg [31:0] _RAND_2022;
  reg [31:0] _RAND_2023;
  reg [31:0] _RAND_2024;
  reg [31:0] _RAND_2025;
  reg [31:0] _RAND_2026;
  reg [31:0] _RAND_2027;
  reg [31:0] _RAND_2028;
  reg [31:0] _RAND_2029;
  reg [31:0] _RAND_2030;
  reg [31:0] _RAND_2031;
  reg [31:0] _RAND_2032;
  reg [31:0] _RAND_2033;
  reg [31:0] _RAND_2034;
  reg [31:0] _RAND_2035;
  reg [31:0] _RAND_2036;
  reg [31:0] _RAND_2037;
  reg [31:0] _RAND_2038;
  reg [31:0] _RAND_2039;
  reg [31:0] _RAND_2040;
  reg [31:0] _RAND_2041;
  reg [31:0] _RAND_2042;
  reg [31:0] _RAND_2043;
  reg [31:0] _RAND_2044;
  reg [31:0] _RAND_2045;
  reg [31:0] _RAND_2046;
  reg [31:0] _RAND_2047;
  reg [31:0] _RAND_2048;
  reg [31:0] _RAND_2049;
  reg [31:0] _RAND_2050;
  reg [31:0] _RAND_2051;
  reg [31:0] _RAND_2052;
  reg [31:0] _RAND_2053;
  reg [31:0] _RAND_2054;
  reg [31:0] _RAND_2055;
  reg [31:0] _RAND_2056;
  reg [31:0] _RAND_2057;
  reg [31:0] _RAND_2058;
  reg [31:0] _RAND_2059;
  reg [31:0] _RAND_2060;
  reg [31:0] _RAND_2061;
  reg [31:0] _RAND_2062;
  reg [31:0] _RAND_2063;
  reg [31:0] _RAND_2064;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] zeroAccumulators_0; // @[BufferAMSNew.scala 14:33]
  reg [7:0] zeroAccumulators_1; // @[BufferAMSNew.scala 14:33]
  reg [7:0] zeroAccumulators_2; // @[BufferAMSNew.scala 14:33]
  reg [7:0] zeroAccumulators_3; // @[BufferAMSNew.scala 14:33]
  reg [7:0] zeroAccumulators_4; // @[BufferAMSNew.scala 14:33]
  reg [7:0] zeroAccumulators_5; // @[BufferAMSNew.scala 14:33]
  reg [7:0] zeroAccumulators_6; // @[BufferAMSNew.scala 14:33]
  reg [7:0] zeroAccumulators_7; // @[BufferAMSNew.scala 14:33]
  reg [3:0] indexAccumulators_0; // @[BufferAMSNew.scala 17:34]
  reg [3:0] indexAccumulators_1; // @[BufferAMSNew.scala 17:34]
  reg [3:0] indexAccumulators_2; // @[BufferAMSNew.scala 17:34]
  reg [3:0] indexAccumulators_3; // @[BufferAMSNew.scala 17:34]
  reg [3:0] indexAccumulators_4; // @[BufferAMSNew.scala 17:34]
  reg [3:0] indexAccumulators_5; // @[BufferAMSNew.scala 17:34]
  reg [3:0] indexAccumulators_6; // @[BufferAMSNew.scala 17:34]
  reg [3:0] indexAccumulators_7; // @[BufferAMSNew.scala 17:34]
  reg [7:0] frameBuffer_0_0; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_1; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_2; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_3; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_4; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_5; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_6; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_7; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_8; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_9; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_10; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_11; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_12; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_13; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_14; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_15; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_16; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_17; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_18; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_19; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_20; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_21; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_22; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_23; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_24; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_25; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_26; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_27; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_28; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_29; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_30; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_31; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_32; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_33; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_34; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_35; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_36; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_37; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_38; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_39; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_40; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_41; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_42; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_43; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_44; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_45; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_46; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_47; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_48; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_49; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_50; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_51; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_52; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_53; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_54; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_55; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_56; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_57; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_58; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_59; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_60; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_61; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_62; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_63; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_64; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_65; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_66; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_67; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_68; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_69; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_70; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_71; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_72; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_73; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_74; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_75; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_76; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_77; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_78; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_79; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_80; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_81; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_82; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_83; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_84; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_85; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_86; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_87; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_88; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_89; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_90; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_91; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_92; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_93; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_94; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_95; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_96; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_97; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_98; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_99; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_100; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_101; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_102; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_103; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_104; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_105; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_106; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_107; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_108; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_109; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_110; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_111; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_112; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_113; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_114; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_115; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_116; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_117; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_118; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_119; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_120; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_121; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_122; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_123; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_124; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_125; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_126; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_0_127; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_0; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_1; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_2; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_3; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_4; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_5; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_6; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_7; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_8; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_9; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_10; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_11; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_12; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_13; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_14; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_15; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_16; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_17; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_18; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_19; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_20; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_21; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_22; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_23; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_24; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_25; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_26; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_27; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_28; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_29; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_30; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_31; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_32; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_33; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_34; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_35; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_36; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_37; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_38; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_39; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_40; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_41; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_42; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_43; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_44; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_45; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_46; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_47; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_48; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_49; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_50; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_51; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_52; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_53; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_54; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_55; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_56; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_57; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_58; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_59; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_60; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_61; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_62; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_63; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_64; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_65; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_66; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_67; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_68; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_69; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_70; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_71; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_72; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_73; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_74; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_75; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_76; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_77; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_78; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_79; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_80; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_81; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_82; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_83; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_84; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_85; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_86; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_87; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_88; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_89; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_90; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_91; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_92; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_93; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_94; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_95; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_96; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_97; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_98; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_99; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_100; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_101; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_102; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_103; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_104; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_105; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_106; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_107; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_108; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_109; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_110; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_111; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_112; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_113; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_114; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_115; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_116; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_117; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_118; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_119; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_120; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_121; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_122; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_123; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_124; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_125; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_126; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_1_127; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_0; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_1; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_2; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_3; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_4; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_5; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_6; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_7; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_8; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_9; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_10; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_11; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_12; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_13; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_14; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_15; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_16; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_17; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_18; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_19; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_20; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_21; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_22; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_23; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_24; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_25; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_26; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_27; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_28; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_29; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_30; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_31; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_32; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_33; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_34; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_35; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_36; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_37; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_38; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_39; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_40; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_41; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_42; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_43; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_44; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_45; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_46; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_47; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_48; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_49; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_50; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_51; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_52; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_53; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_54; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_55; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_56; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_57; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_58; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_59; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_60; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_61; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_62; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_63; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_64; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_65; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_66; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_67; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_68; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_69; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_70; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_71; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_72; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_73; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_74; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_75; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_76; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_77; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_78; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_79; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_80; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_81; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_82; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_83; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_84; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_85; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_86; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_87; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_88; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_89; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_90; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_91; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_92; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_93; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_94; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_95; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_96; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_97; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_98; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_99; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_100; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_101; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_102; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_103; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_104; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_105; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_106; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_107; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_108; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_109; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_110; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_111; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_112; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_113; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_114; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_115; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_116; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_117; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_118; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_119; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_120; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_121; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_122; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_123; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_124; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_125; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_126; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_2_127; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_0; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_1; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_2; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_3; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_4; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_5; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_6; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_7; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_8; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_9; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_10; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_11; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_12; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_13; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_14; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_15; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_16; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_17; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_18; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_19; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_20; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_21; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_22; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_23; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_24; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_25; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_26; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_27; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_28; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_29; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_30; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_31; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_32; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_33; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_34; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_35; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_36; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_37; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_38; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_39; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_40; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_41; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_42; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_43; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_44; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_45; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_46; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_47; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_48; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_49; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_50; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_51; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_52; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_53; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_54; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_55; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_56; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_57; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_58; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_59; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_60; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_61; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_62; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_63; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_64; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_65; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_66; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_67; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_68; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_69; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_70; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_71; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_72; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_73; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_74; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_75; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_76; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_77; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_78; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_79; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_80; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_81; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_82; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_83; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_84; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_85; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_86; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_87; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_88; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_89; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_90; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_91; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_92; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_93; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_94; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_95; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_96; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_97; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_98; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_99; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_100; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_101; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_102; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_103; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_104; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_105; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_106; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_107; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_108; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_109; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_110; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_111; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_112; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_113; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_114; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_115; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_116; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_117; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_118; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_119; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_120; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_121; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_122; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_123; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_124; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_125; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_126; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_3_127; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_0; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_1; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_2; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_3; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_4; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_5; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_6; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_7; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_8; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_9; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_10; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_11; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_12; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_13; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_14; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_15; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_16; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_17; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_18; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_19; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_20; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_21; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_22; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_23; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_24; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_25; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_26; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_27; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_28; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_29; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_30; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_31; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_32; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_33; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_34; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_35; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_36; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_37; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_38; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_39; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_40; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_41; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_42; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_43; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_44; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_45; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_46; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_47; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_48; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_49; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_50; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_51; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_52; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_53; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_54; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_55; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_56; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_57; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_58; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_59; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_60; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_61; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_62; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_63; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_64; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_65; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_66; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_67; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_68; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_69; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_70; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_71; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_72; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_73; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_74; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_75; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_76; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_77; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_78; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_79; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_80; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_81; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_82; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_83; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_84; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_85; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_86; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_87; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_88; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_89; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_90; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_91; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_92; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_93; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_94; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_95; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_96; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_97; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_98; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_99; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_100; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_101; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_102; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_103; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_104; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_105; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_106; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_107; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_108; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_109; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_110; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_111; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_112; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_113; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_114; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_115; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_116; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_117; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_118; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_119; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_120; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_121; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_122; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_123; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_124; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_125; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_126; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_4_127; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_0; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_1; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_2; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_3; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_4; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_5; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_6; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_7; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_8; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_9; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_10; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_11; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_12; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_13; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_14; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_15; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_16; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_17; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_18; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_19; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_20; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_21; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_22; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_23; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_24; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_25; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_26; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_27; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_28; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_29; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_30; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_31; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_32; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_33; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_34; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_35; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_36; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_37; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_38; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_39; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_40; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_41; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_42; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_43; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_44; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_45; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_46; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_47; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_48; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_49; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_50; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_51; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_52; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_53; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_54; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_55; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_56; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_57; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_58; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_59; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_60; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_61; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_62; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_63; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_64; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_65; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_66; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_67; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_68; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_69; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_70; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_71; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_72; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_73; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_74; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_75; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_76; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_77; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_78; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_79; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_80; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_81; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_82; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_83; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_84; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_85; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_86; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_87; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_88; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_89; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_90; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_91; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_92; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_93; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_94; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_95; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_96; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_97; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_98; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_99; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_100; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_101; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_102; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_103; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_104; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_105; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_106; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_107; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_108; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_109; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_110; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_111; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_112; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_113; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_114; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_115; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_116; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_117; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_118; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_119; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_120; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_121; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_122; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_123; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_124; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_125; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_126; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_5_127; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_0; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_1; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_2; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_3; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_4; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_5; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_6; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_7; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_8; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_9; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_10; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_11; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_12; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_13; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_14; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_15; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_16; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_17; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_18; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_19; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_20; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_21; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_22; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_23; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_24; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_25; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_26; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_27; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_28; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_29; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_30; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_31; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_32; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_33; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_34; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_35; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_36; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_37; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_38; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_39; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_40; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_41; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_42; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_43; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_44; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_45; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_46; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_47; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_48; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_49; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_50; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_51; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_52; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_53; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_54; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_55; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_56; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_57; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_58; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_59; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_60; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_61; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_62; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_63; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_64; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_65; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_66; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_67; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_68; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_69; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_70; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_71; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_72; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_73; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_74; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_75; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_76; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_77; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_78; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_79; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_80; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_81; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_82; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_83; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_84; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_85; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_86; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_87; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_88; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_89; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_90; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_91; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_92; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_93; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_94; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_95; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_96; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_97; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_98; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_99; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_100; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_101; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_102; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_103; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_104; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_105; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_106; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_107; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_108; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_109; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_110; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_111; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_112; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_113; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_114; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_115; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_116; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_117; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_118; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_119; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_120; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_121; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_122; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_123; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_124; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_125; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_126; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_6_127; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_0; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_1; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_2; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_3; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_4; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_5; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_6; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_7; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_8; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_9; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_10; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_11; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_12; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_13; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_14; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_15; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_16; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_17; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_18; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_19; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_20; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_21; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_22; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_23; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_24; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_25; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_26; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_27; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_28; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_29; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_30; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_31; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_32; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_33; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_34; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_35; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_36; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_37; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_38; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_39; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_40; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_41; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_42; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_43; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_44; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_45; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_46; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_47; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_48; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_49; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_50; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_51; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_52; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_53; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_54; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_55; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_56; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_57; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_58; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_59; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_60; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_61; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_62; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_63; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_64; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_65; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_66; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_67; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_68; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_69; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_70; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_71; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_72; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_73; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_74; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_75; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_76; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_77; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_78; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_79; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_80; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_81; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_82; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_83; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_84; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_85; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_86; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_87; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_88; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_89; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_90; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_91; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_92; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_93; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_94; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_95; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_96; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_97; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_98; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_99; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_100; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_101; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_102; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_103; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_104; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_105; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_106; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_107; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_108; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_109; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_110; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_111; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_112; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_113; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_114; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_115; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_116; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_117; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_118; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_119; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_120; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_121; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_122; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_123; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_124; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_125; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_126; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_7_127; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_0; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_1; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_2; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_3; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_4; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_5; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_6; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_7; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_8; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_9; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_10; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_11; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_12; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_13; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_14; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_15; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_16; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_17; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_18; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_19; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_20; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_21; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_22; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_23; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_24; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_25; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_26; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_27; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_28; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_29; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_30; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_31; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_32; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_33; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_34; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_35; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_36; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_37; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_38; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_39; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_40; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_41; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_42; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_43; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_44; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_45; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_46; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_47; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_48; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_49; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_50; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_51; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_52; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_53; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_54; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_55; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_56; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_57; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_58; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_59; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_60; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_61; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_62; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_63; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_64; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_65; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_66; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_67; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_68; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_69; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_70; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_71; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_72; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_73; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_74; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_75; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_76; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_77; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_78; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_79; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_80; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_81; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_82; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_83; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_84; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_85; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_86; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_87; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_88; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_89; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_90; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_91; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_92; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_93; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_94; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_95; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_96; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_97; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_98; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_99; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_100; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_101; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_102; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_103; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_104; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_105; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_106; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_107; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_108; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_109; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_110; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_111; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_112; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_113; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_114; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_115; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_116; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_117; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_118; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_119; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_120; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_121; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_122; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_123; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_124; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_125; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_126; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_8_127; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_0; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_1; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_2; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_3; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_4; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_5; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_6; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_7; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_8; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_9; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_10; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_11; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_12; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_13; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_14; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_15; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_16; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_17; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_18; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_19; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_20; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_21; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_22; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_23; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_24; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_25; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_26; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_27; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_28; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_29; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_30; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_31; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_32; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_33; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_34; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_35; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_36; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_37; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_38; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_39; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_40; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_41; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_42; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_43; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_44; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_45; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_46; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_47; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_48; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_49; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_50; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_51; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_52; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_53; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_54; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_55; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_56; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_57; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_58; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_59; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_60; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_61; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_62; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_63; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_64; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_65; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_66; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_67; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_68; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_69; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_70; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_71; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_72; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_73; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_74; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_75; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_76; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_77; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_78; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_79; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_80; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_81; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_82; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_83; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_84; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_85; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_86; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_87; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_88; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_89; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_90; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_91; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_92; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_93; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_94; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_95; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_96; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_97; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_98; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_99; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_100; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_101; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_102; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_103; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_104; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_105; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_106; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_107; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_108; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_109; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_110; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_111; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_112; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_113; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_114; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_115; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_116; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_117; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_118; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_119; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_120; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_121; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_122; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_123; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_124; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_125; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_126; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_9_127; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_0; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_1; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_2; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_3; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_4; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_5; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_6; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_7; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_8; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_9; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_10; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_11; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_12; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_13; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_14; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_15; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_16; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_17; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_18; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_19; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_20; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_21; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_22; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_23; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_24; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_25; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_26; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_27; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_28; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_29; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_30; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_31; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_32; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_33; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_34; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_35; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_36; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_37; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_38; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_39; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_40; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_41; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_42; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_43; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_44; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_45; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_46; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_47; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_48; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_49; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_50; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_51; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_52; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_53; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_54; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_55; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_56; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_57; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_58; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_59; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_60; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_61; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_62; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_63; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_64; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_65; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_66; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_67; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_68; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_69; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_70; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_71; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_72; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_73; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_74; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_75; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_76; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_77; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_78; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_79; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_80; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_81; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_82; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_83; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_84; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_85; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_86; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_87; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_88; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_89; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_90; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_91; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_92; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_93; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_94; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_95; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_96; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_97; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_98; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_99; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_100; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_101; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_102; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_103; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_104; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_105; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_106; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_107; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_108; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_109; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_110; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_111; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_112; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_113; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_114; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_115; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_116; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_117; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_118; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_119; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_120; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_121; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_122; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_123; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_124; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_125; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_126; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_10_127; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_0; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_1; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_2; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_3; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_4; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_5; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_6; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_7; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_8; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_9; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_10; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_11; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_12; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_13; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_14; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_15; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_16; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_17; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_18; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_19; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_20; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_21; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_22; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_23; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_24; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_25; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_26; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_27; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_28; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_29; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_30; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_31; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_32; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_33; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_34; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_35; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_36; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_37; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_38; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_39; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_40; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_41; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_42; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_43; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_44; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_45; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_46; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_47; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_48; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_49; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_50; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_51; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_52; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_53; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_54; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_55; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_56; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_57; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_58; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_59; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_60; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_61; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_62; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_63; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_64; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_65; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_66; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_67; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_68; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_69; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_70; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_71; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_72; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_73; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_74; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_75; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_76; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_77; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_78; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_79; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_80; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_81; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_82; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_83; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_84; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_85; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_86; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_87; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_88; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_89; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_90; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_91; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_92; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_93; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_94; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_95; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_96; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_97; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_98; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_99; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_100; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_101; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_102; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_103; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_104; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_105; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_106; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_107; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_108; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_109; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_110; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_111; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_112; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_113; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_114; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_115; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_116; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_117; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_118; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_119; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_120; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_121; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_122; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_123; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_124; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_125; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_126; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_11_127; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_0; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_1; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_2; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_3; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_4; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_5; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_6; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_7; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_8; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_9; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_10; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_11; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_12; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_13; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_14; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_15; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_16; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_17; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_18; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_19; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_20; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_21; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_22; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_23; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_24; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_25; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_26; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_27; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_28; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_29; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_30; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_31; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_32; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_33; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_34; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_35; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_36; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_37; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_38; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_39; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_40; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_41; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_42; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_43; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_44; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_45; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_46; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_47; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_48; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_49; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_50; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_51; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_52; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_53; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_54; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_55; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_56; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_57; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_58; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_59; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_60; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_61; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_62; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_63; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_64; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_65; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_66; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_67; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_68; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_69; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_70; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_71; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_72; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_73; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_74; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_75; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_76; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_77; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_78; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_79; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_80; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_81; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_82; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_83; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_84; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_85; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_86; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_87; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_88; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_89; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_90; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_91; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_92; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_93; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_94; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_95; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_96; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_97; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_98; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_99; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_100; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_101; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_102; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_103; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_104; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_105; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_106; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_107; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_108; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_109; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_110; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_111; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_112; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_113; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_114; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_115; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_116; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_117; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_118; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_119; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_120; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_121; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_122; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_123; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_124; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_125; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_126; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_12_127; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_0; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_1; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_2; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_3; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_4; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_5; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_6; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_7; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_8; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_9; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_10; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_11; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_12; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_13; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_14; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_15; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_16; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_17; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_18; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_19; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_20; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_21; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_22; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_23; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_24; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_25; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_26; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_27; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_28; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_29; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_30; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_31; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_32; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_33; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_34; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_35; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_36; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_37; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_38; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_39; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_40; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_41; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_42; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_43; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_44; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_45; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_46; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_47; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_48; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_49; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_50; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_51; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_52; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_53; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_54; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_55; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_56; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_57; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_58; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_59; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_60; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_61; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_62; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_63; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_64; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_65; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_66; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_67; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_68; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_69; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_70; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_71; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_72; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_73; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_74; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_75; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_76; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_77; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_78; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_79; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_80; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_81; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_82; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_83; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_84; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_85; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_86; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_87; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_88; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_89; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_90; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_91; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_92; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_93; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_94; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_95; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_96; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_97; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_98; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_99; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_100; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_101; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_102; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_103; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_104; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_105; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_106; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_107; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_108; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_109; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_110; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_111; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_112; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_113; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_114; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_115; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_116; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_117; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_118; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_119; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_120; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_121; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_122; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_123; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_124; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_125; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_126; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_13_127; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_0; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_1; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_2; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_3; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_4; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_5; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_6; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_7; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_8; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_9; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_10; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_11; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_12; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_13; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_14; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_15; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_16; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_17; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_18; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_19; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_20; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_21; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_22; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_23; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_24; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_25; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_26; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_27; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_28; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_29; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_30; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_31; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_32; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_33; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_34; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_35; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_36; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_37; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_38; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_39; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_40; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_41; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_42; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_43; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_44; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_45; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_46; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_47; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_48; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_49; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_50; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_51; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_52; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_53; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_54; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_55; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_56; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_57; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_58; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_59; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_60; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_61; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_62; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_63; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_64; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_65; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_66; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_67; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_68; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_69; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_70; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_71; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_72; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_73; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_74; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_75; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_76; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_77; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_78; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_79; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_80; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_81; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_82; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_83; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_84; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_85; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_86; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_87; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_88; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_89; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_90; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_91; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_92; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_93; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_94; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_95; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_96; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_97; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_98; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_99; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_100; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_101; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_102; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_103; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_104; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_105; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_106; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_107; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_108; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_109; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_110; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_111; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_112; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_113; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_114; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_115; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_116; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_117; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_118; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_119; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_120; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_121; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_122; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_123; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_124; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_125; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_126; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_14_127; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_0; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_1; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_2; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_3; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_4; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_5; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_6; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_7; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_8; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_9; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_10; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_11; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_12; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_13; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_14; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_15; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_16; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_17; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_18; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_19; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_20; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_21; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_22; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_23; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_24; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_25; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_26; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_27; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_28; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_29; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_30; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_31; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_32; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_33; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_34; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_35; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_36; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_37; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_38; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_39; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_40; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_41; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_42; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_43; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_44; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_45; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_46; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_47; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_48; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_49; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_50; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_51; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_52; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_53; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_54; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_55; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_56; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_57; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_58; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_59; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_60; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_61; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_62; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_63; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_64; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_65; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_66; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_67; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_68; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_69; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_70; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_71; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_72; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_73; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_74; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_75; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_76; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_77; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_78; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_79; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_80; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_81; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_82; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_83; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_84; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_85; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_86; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_87; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_88; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_89; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_90; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_91; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_92; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_93; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_94; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_95; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_96; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_97; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_98; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_99; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_100; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_101; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_102; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_103; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_104; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_105; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_106; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_107; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_108; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_109; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_110; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_111; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_112; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_113; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_114; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_115; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_116; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_117; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_118; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_119; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_120; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_121; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_122; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_123; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_124; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_125; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_126; // @[BufferAMSNew.scala 20:24]
  reg [7:0] frameBuffer_15_127; // @[BufferAMSNew.scala 20:24]
  reg [3:0] lineCounter; // @[BufferAMSNew.scala 21:28]
  wire [3:0] _lineCounter_T_1 = lineCounter + 4'h1; // @[BufferAMSNew.scala 33:32]
  wire [1:0] _zeroCount_T_16 = {{1'd0}, io_adcValues_0 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [1:0] _GEN_4225 = {{1'd0}, io_adcValues_1 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [2:0] _zeroCount_T_17 = _zeroCount_T_16 + _GEN_4225; // @[BufferAMSNew.scala 38:70]
  wire [2:0] _GEN_4226 = {{2'd0}, io_adcValues_2 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [3:0] _zeroCount_T_18 = _zeroCount_T_17 + _GEN_4226; // @[BufferAMSNew.scala 38:70]
  wire [3:0] _GEN_4227 = {{3'd0}, io_adcValues_3 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [4:0] _zeroCount_T_19 = _zeroCount_T_18 + _GEN_4227; // @[BufferAMSNew.scala 38:70]
  wire [4:0] _GEN_4228 = {{4'd0}, io_adcValues_4 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [5:0] _zeroCount_T_20 = _zeroCount_T_19 + _GEN_4228; // @[BufferAMSNew.scala 38:70]
  wire [5:0] _GEN_4229 = {{5'd0}, io_adcValues_5 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [6:0] _zeroCount_T_21 = _zeroCount_T_20 + _GEN_4229; // @[BufferAMSNew.scala 38:70]
  wire [6:0] _GEN_4230 = {{6'd0}, io_adcValues_6 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [7:0] _zeroCount_T_22 = _zeroCount_T_21 + _GEN_4230; // @[BufferAMSNew.scala 38:70]
  wire [7:0] _GEN_4231 = {{7'd0}, io_adcValues_7 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [8:0] _zeroCount_T_23 = _zeroCount_T_22 + _GEN_4231; // @[BufferAMSNew.scala 38:70]
  wire [8:0] _GEN_4232 = {{8'd0}, io_adcValues_8 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [9:0] _zeroCount_T_24 = _zeroCount_T_23 + _GEN_4232; // @[BufferAMSNew.scala 38:70]
  wire [9:0] _GEN_4233 = {{9'd0}, io_adcValues_9 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [10:0] _zeroCount_T_25 = _zeroCount_T_24 + _GEN_4233; // @[BufferAMSNew.scala 38:70]
  wire [10:0] _GEN_4234 = {{10'd0}, io_adcValues_10 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [11:0] _zeroCount_T_26 = _zeroCount_T_25 + _GEN_4234; // @[BufferAMSNew.scala 38:70]
  wire [11:0] _GEN_4235 = {{11'd0}, io_adcValues_11 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [12:0] _zeroCount_T_27 = _zeroCount_T_26 + _GEN_4235; // @[BufferAMSNew.scala 38:70]
  wire [12:0] _GEN_4236 = {{12'd0}, io_adcValues_12 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [13:0] _zeroCount_T_28 = _zeroCount_T_27 + _GEN_4236; // @[BufferAMSNew.scala 38:70]
  wire [13:0] _GEN_4237 = {{13'd0}, io_adcValues_13 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [14:0] _zeroCount_T_29 = _zeroCount_T_28 + _GEN_4237; // @[BufferAMSNew.scala 38:70]
  wire [14:0] _GEN_4238 = {{14'd0}, io_adcValues_14 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [15:0] _zeroCount_T_30 = _zeroCount_T_29 + _GEN_4238; // @[BufferAMSNew.scala 38:70]
  wire [15:0] _GEN_4239 = {{15'd0}, io_adcValues_15 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [16:0] zeroCount = _zeroCount_T_30 + _GEN_4239; // @[BufferAMSNew.scala 38:70]
  wire [16:0] _GEN_4240 = {{9'd0}, zeroAccumulators_0}; // @[BufferAMSNew.scala 41:50]
  wire [16:0] _zeroAccumulators_0_T_1 = _GEN_4240 + zeroCount; // @[BufferAMSNew.scala 41:50]
  wire [1:0] _zeroCount_T_47 = {{1'd0}, io_adcValues_16 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [1:0] _GEN_4241 = {{1'd0}, io_adcValues_17 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [2:0] _zeroCount_T_48 = _zeroCount_T_47 + _GEN_4241; // @[BufferAMSNew.scala 38:70]
  wire [2:0] _GEN_4242 = {{2'd0}, io_adcValues_18 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [3:0] _zeroCount_T_49 = _zeroCount_T_48 + _GEN_4242; // @[BufferAMSNew.scala 38:70]
  wire [3:0] _GEN_4243 = {{3'd0}, io_adcValues_19 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [4:0] _zeroCount_T_50 = _zeroCount_T_49 + _GEN_4243; // @[BufferAMSNew.scala 38:70]
  wire [4:0] _GEN_4244 = {{4'd0}, io_adcValues_20 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [5:0] _zeroCount_T_51 = _zeroCount_T_50 + _GEN_4244; // @[BufferAMSNew.scala 38:70]
  wire [5:0] _GEN_4245 = {{5'd0}, io_adcValues_21 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [6:0] _zeroCount_T_52 = _zeroCount_T_51 + _GEN_4245; // @[BufferAMSNew.scala 38:70]
  wire [6:0] _GEN_4246 = {{6'd0}, io_adcValues_22 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [7:0] _zeroCount_T_53 = _zeroCount_T_52 + _GEN_4246; // @[BufferAMSNew.scala 38:70]
  wire [7:0] _GEN_4247 = {{7'd0}, io_adcValues_23 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [8:0] _zeroCount_T_54 = _zeroCount_T_53 + _GEN_4247; // @[BufferAMSNew.scala 38:70]
  wire [8:0] _GEN_4248 = {{8'd0}, io_adcValues_24 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [9:0] _zeroCount_T_55 = _zeroCount_T_54 + _GEN_4248; // @[BufferAMSNew.scala 38:70]
  wire [9:0] _GEN_4249 = {{9'd0}, io_adcValues_25 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [10:0] _zeroCount_T_56 = _zeroCount_T_55 + _GEN_4249; // @[BufferAMSNew.scala 38:70]
  wire [10:0] _GEN_4250 = {{10'd0}, io_adcValues_26 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [11:0] _zeroCount_T_57 = _zeroCount_T_56 + _GEN_4250; // @[BufferAMSNew.scala 38:70]
  wire [11:0] _GEN_4251 = {{11'd0}, io_adcValues_27 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [12:0] _zeroCount_T_58 = _zeroCount_T_57 + _GEN_4251; // @[BufferAMSNew.scala 38:70]
  wire [12:0] _GEN_4252 = {{12'd0}, io_adcValues_28 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [13:0] _zeroCount_T_59 = _zeroCount_T_58 + _GEN_4252; // @[BufferAMSNew.scala 38:70]
  wire [13:0] _GEN_4253 = {{13'd0}, io_adcValues_29 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [14:0] _zeroCount_T_60 = _zeroCount_T_59 + _GEN_4253; // @[BufferAMSNew.scala 38:70]
  wire [14:0] _GEN_4254 = {{14'd0}, io_adcValues_30 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [15:0] _zeroCount_T_61 = _zeroCount_T_60 + _GEN_4254; // @[BufferAMSNew.scala 38:70]
  wire [15:0] _GEN_4255 = {{15'd0}, io_adcValues_31 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [16:0] zeroCount_1 = _zeroCount_T_61 + _GEN_4255; // @[BufferAMSNew.scala 38:70]
  wire [16:0] _GEN_4256 = {{9'd0}, zeroAccumulators_1}; // @[BufferAMSNew.scala 41:50]
  wire [16:0] _zeroAccumulators_1_T_1 = _GEN_4256 + zeroCount_1; // @[BufferAMSNew.scala 41:50]
  wire [1:0] _zeroCount_T_78 = {{1'd0}, io_adcValues_32 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [1:0] _GEN_4257 = {{1'd0}, io_adcValues_33 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [2:0] _zeroCount_T_79 = _zeroCount_T_78 + _GEN_4257; // @[BufferAMSNew.scala 38:70]
  wire [2:0] _GEN_4258 = {{2'd0}, io_adcValues_34 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [3:0] _zeroCount_T_80 = _zeroCount_T_79 + _GEN_4258; // @[BufferAMSNew.scala 38:70]
  wire [3:0] _GEN_4259 = {{3'd0}, io_adcValues_35 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [4:0] _zeroCount_T_81 = _zeroCount_T_80 + _GEN_4259; // @[BufferAMSNew.scala 38:70]
  wire [4:0] _GEN_4260 = {{4'd0}, io_adcValues_36 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [5:0] _zeroCount_T_82 = _zeroCount_T_81 + _GEN_4260; // @[BufferAMSNew.scala 38:70]
  wire [5:0] _GEN_4261 = {{5'd0}, io_adcValues_37 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [6:0] _zeroCount_T_83 = _zeroCount_T_82 + _GEN_4261; // @[BufferAMSNew.scala 38:70]
  wire [6:0] _GEN_4262 = {{6'd0}, io_adcValues_38 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [7:0] _zeroCount_T_84 = _zeroCount_T_83 + _GEN_4262; // @[BufferAMSNew.scala 38:70]
  wire [7:0] _GEN_4263 = {{7'd0}, io_adcValues_39 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [8:0] _zeroCount_T_85 = _zeroCount_T_84 + _GEN_4263; // @[BufferAMSNew.scala 38:70]
  wire [8:0] _GEN_4264 = {{8'd0}, io_adcValues_40 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [9:0] _zeroCount_T_86 = _zeroCount_T_85 + _GEN_4264; // @[BufferAMSNew.scala 38:70]
  wire [9:0] _GEN_4265 = {{9'd0}, io_adcValues_41 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [10:0] _zeroCount_T_87 = _zeroCount_T_86 + _GEN_4265; // @[BufferAMSNew.scala 38:70]
  wire [10:0] _GEN_4266 = {{10'd0}, io_adcValues_42 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [11:0] _zeroCount_T_88 = _zeroCount_T_87 + _GEN_4266; // @[BufferAMSNew.scala 38:70]
  wire [11:0] _GEN_4267 = {{11'd0}, io_adcValues_43 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [12:0] _zeroCount_T_89 = _zeroCount_T_88 + _GEN_4267; // @[BufferAMSNew.scala 38:70]
  wire [12:0] _GEN_4268 = {{12'd0}, io_adcValues_44 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [13:0] _zeroCount_T_90 = _zeroCount_T_89 + _GEN_4268; // @[BufferAMSNew.scala 38:70]
  wire [13:0] _GEN_4269 = {{13'd0}, io_adcValues_45 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [14:0] _zeroCount_T_91 = _zeroCount_T_90 + _GEN_4269; // @[BufferAMSNew.scala 38:70]
  wire [14:0] _GEN_4270 = {{14'd0}, io_adcValues_46 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [15:0] _zeroCount_T_92 = _zeroCount_T_91 + _GEN_4270; // @[BufferAMSNew.scala 38:70]
  wire [15:0] _GEN_4271 = {{15'd0}, io_adcValues_47 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [16:0] zeroCount_2 = _zeroCount_T_92 + _GEN_4271; // @[BufferAMSNew.scala 38:70]
  wire [16:0] _GEN_4272 = {{9'd0}, zeroAccumulators_2}; // @[BufferAMSNew.scala 41:50]
  wire [16:0] _zeroAccumulators_2_T_1 = _GEN_4272 + zeroCount_2; // @[BufferAMSNew.scala 41:50]
  wire [1:0] _zeroCount_T_109 = {{1'd0}, io_adcValues_48 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [1:0] _GEN_4273 = {{1'd0}, io_adcValues_49 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [2:0] _zeroCount_T_110 = _zeroCount_T_109 + _GEN_4273; // @[BufferAMSNew.scala 38:70]
  wire [2:0] _GEN_4274 = {{2'd0}, io_adcValues_50 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [3:0] _zeroCount_T_111 = _zeroCount_T_110 + _GEN_4274; // @[BufferAMSNew.scala 38:70]
  wire [3:0] _GEN_4275 = {{3'd0}, io_adcValues_51 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [4:0] _zeroCount_T_112 = _zeroCount_T_111 + _GEN_4275; // @[BufferAMSNew.scala 38:70]
  wire [4:0] _GEN_4276 = {{4'd0}, io_adcValues_52 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [5:0] _zeroCount_T_113 = _zeroCount_T_112 + _GEN_4276; // @[BufferAMSNew.scala 38:70]
  wire [5:0] _GEN_4277 = {{5'd0}, io_adcValues_53 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [6:0] _zeroCount_T_114 = _zeroCount_T_113 + _GEN_4277; // @[BufferAMSNew.scala 38:70]
  wire [6:0] _GEN_4278 = {{6'd0}, io_adcValues_54 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [7:0] _zeroCount_T_115 = _zeroCount_T_114 + _GEN_4278; // @[BufferAMSNew.scala 38:70]
  wire [7:0] _GEN_4279 = {{7'd0}, io_adcValues_55 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [8:0] _zeroCount_T_116 = _zeroCount_T_115 + _GEN_4279; // @[BufferAMSNew.scala 38:70]
  wire [8:0] _GEN_4280 = {{8'd0}, io_adcValues_56 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [9:0] _zeroCount_T_117 = _zeroCount_T_116 + _GEN_4280; // @[BufferAMSNew.scala 38:70]
  wire [9:0] _GEN_4281 = {{9'd0}, io_adcValues_57 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [10:0] _zeroCount_T_118 = _zeroCount_T_117 + _GEN_4281; // @[BufferAMSNew.scala 38:70]
  wire [10:0] _GEN_4282 = {{10'd0}, io_adcValues_58 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [11:0] _zeroCount_T_119 = _zeroCount_T_118 + _GEN_4282; // @[BufferAMSNew.scala 38:70]
  wire [11:0] _GEN_4283 = {{11'd0}, io_adcValues_59 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [12:0] _zeroCount_T_120 = _zeroCount_T_119 + _GEN_4283; // @[BufferAMSNew.scala 38:70]
  wire [12:0] _GEN_4284 = {{12'd0}, io_adcValues_60 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [13:0] _zeroCount_T_121 = _zeroCount_T_120 + _GEN_4284; // @[BufferAMSNew.scala 38:70]
  wire [13:0] _GEN_4285 = {{13'd0}, io_adcValues_61 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [14:0] _zeroCount_T_122 = _zeroCount_T_121 + _GEN_4285; // @[BufferAMSNew.scala 38:70]
  wire [14:0] _GEN_4286 = {{14'd0}, io_adcValues_62 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [15:0] _zeroCount_T_123 = _zeroCount_T_122 + _GEN_4286; // @[BufferAMSNew.scala 38:70]
  wire [15:0] _GEN_4287 = {{15'd0}, io_adcValues_63 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [16:0] zeroCount_3 = _zeroCount_T_123 + _GEN_4287; // @[BufferAMSNew.scala 38:70]
  wire [16:0] _GEN_4288 = {{9'd0}, zeroAccumulators_3}; // @[BufferAMSNew.scala 41:50]
  wire [16:0] _zeroAccumulators_3_T_1 = _GEN_4288 + zeroCount_3; // @[BufferAMSNew.scala 41:50]
  wire [1:0] _zeroCount_T_140 = {{1'd0}, io_adcValues_64 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [1:0] _GEN_4289 = {{1'd0}, io_adcValues_65 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [2:0] _zeroCount_T_141 = _zeroCount_T_140 + _GEN_4289; // @[BufferAMSNew.scala 38:70]
  wire [2:0] _GEN_4290 = {{2'd0}, io_adcValues_66 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [3:0] _zeroCount_T_142 = _zeroCount_T_141 + _GEN_4290; // @[BufferAMSNew.scala 38:70]
  wire [3:0] _GEN_4291 = {{3'd0}, io_adcValues_67 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [4:0] _zeroCount_T_143 = _zeroCount_T_142 + _GEN_4291; // @[BufferAMSNew.scala 38:70]
  wire [4:0] _GEN_4292 = {{4'd0}, io_adcValues_68 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [5:0] _zeroCount_T_144 = _zeroCount_T_143 + _GEN_4292; // @[BufferAMSNew.scala 38:70]
  wire [5:0] _GEN_4293 = {{5'd0}, io_adcValues_69 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [6:0] _zeroCount_T_145 = _zeroCount_T_144 + _GEN_4293; // @[BufferAMSNew.scala 38:70]
  wire [6:0] _GEN_4294 = {{6'd0}, io_adcValues_70 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [7:0] _zeroCount_T_146 = _zeroCount_T_145 + _GEN_4294; // @[BufferAMSNew.scala 38:70]
  wire [7:0] _GEN_4295 = {{7'd0}, io_adcValues_71 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [8:0] _zeroCount_T_147 = _zeroCount_T_146 + _GEN_4295; // @[BufferAMSNew.scala 38:70]
  wire [8:0] _GEN_4296 = {{8'd0}, io_adcValues_72 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [9:0] _zeroCount_T_148 = _zeroCount_T_147 + _GEN_4296; // @[BufferAMSNew.scala 38:70]
  wire [9:0] _GEN_4297 = {{9'd0}, io_adcValues_73 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [10:0] _zeroCount_T_149 = _zeroCount_T_148 + _GEN_4297; // @[BufferAMSNew.scala 38:70]
  wire [10:0] _GEN_4298 = {{10'd0}, io_adcValues_74 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [11:0] _zeroCount_T_150 = _zeroCount_T_149 + _GEN_4298; // @[BufferAMSNew.scala 38:70]
  wire [11:0] _GEN_4299 = {{11'd0}, io_adcValues_75 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [12:0] _zeroCount_T_151 = _zeroCount_T_150 + _GEN_4299; // @[BufferAMSNew.scala 38:70]
  wire [12:0] _GEN_4300 = {{12'd0}, io_adcValues_76 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [13:0] _zeroCount_T_152 = _zeroCount_T_151 + _GEN_4300; // @[BufferAMSNew.scala 38:70]
  wire [13:0] _GEN_4301 = {{13'd0}, io_adcValues_77 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [14:0] _zeroCount_T_153 = _zeroCount_T_152 + _GEN_4301; // @[BufferAMSNew.scala 38:70]
  wire [14:0] _GEN_4302 = {{14'd0}, io_adcValues_78 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [15:0] _zeroCount_T_154 = _zeroCount_T_153 + _GEN_4302; // @[BufferAMSNew.scala 38:70]
  wire [15:0] _GEN_4303 = {{15'd0}, io_adcValues_79 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [16:0] zeroCount_4 = _zeroCount_T_154 + _GEN_4303; // @[BufferAMSNew.scala 38:70]
  wire [16:0] _GEN_4304 = {{9'd0}, zeroAccumulators_4}; // @[BufferAMSNew.scala 41:50]
  wire [16:0] _zeroAccumulators_4_T_1 = _GEN_4304 + zeroCount_4; // @[BufferAMSNew.scala 41:50]
  wire [1:0] _zeroCount_T_171 = {{1'd0}, io_adcValues_80 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [1:0] _GEN_4305 = {{1'd0}, io_adcValues_81 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [2:0] _zeroCount_T_172 = _zeroCount_T_171 + _GEN_4305; // @[BufferAMSNew.scala 38:70]
  wire [2:0] _GEN_4306 = {{2'd0}, io_adcValues_82 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [3:0] _zeroCount_T_173 = _zeroCount_T_172 + _GEN_4306; // @[BufferAMSNew.scala 38:70]
  wire [3:0] _GEN_4307 = {{3'd0}, io_adcValues_83 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [4:0] _zeroCount_T_174 = _zeroCount_T_173 + _GEN_4307; // @[BufferAMSNew.scala 38:70]
  wire [4:0] _GEN_4308 = {{4'd0}, io_adcValues_84 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [5:0] _zeroCount_T_175 = _zeroCount_T_174 + _GEN_4308; // @[BufferAMSNew.scala 38:70]
  wire [5:0] _GEN_4309 = {{5'd0}, io_adcValues_85 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [6:0] _zeroCount_T_176 = _zeroCount_T_175 + _GEN_4309; // @[BufferAMSNew.scala 38:70]
  wire [6:0] _GEN_4310 = {{6'd0}, io_adcValues_86 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [7:0] _zeroCount_T_177 = _zeroCount_T_176 + _GEN_4310; // @[BufferAMSNew.scala 38:70]
  wire [7:0] _GEN_4311 = {{7'd0}, io_adcValues_87 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [8:0] _zeroCount_T_178 = _zeroCount_T_177 + _GEN_4311; // @[BufferAMSNew.scala 38:70]
  wire [8:0] _GEN_4312 = {{8'd0}, io_adcValues_88 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [9:0] _zeroCount_T_179 = _zeroCount_T_178 + _GEN_4312; // @[BufferAMSNew.scala 38:70]
  wire [9:0] _GEN_4313 = {{9'd0}, io_adcValues_89 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [10:0] _zeroCount_T_180 = _zeroCount_T_179 + _GEN_4313; // @[BufferAMSNew.scala 38:70]
  wire [10:0] _GEN_4314 = {{10'd0}, io_adcValues_90 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [11:0] _zeroCount_T_181 = _zeroCount_T_180 + _GEN_4314; // @[BufferAMSNew.scala 38:70]
  wire [11:0] _GEN_4315 = {{11'd0}, io_adcValues_91 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [12:0] _zeroCount_T_182 = _zeroCount_T_181 + _GEN_4315; // @[BufferAMSNew.scala 38:70]
  wire [12:0] _GEN_4316 = {{12'd0}, io_adcValues_92 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [13:0] _zeroCount_T_183 = _zeroCount_T_182 + _GEN_4316; // @[BufferAMSNew.scala 38:70]
  wire [13:0] _GEN_4317 = {{13'd0}, io_adcValues_93 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [14:0] _zeroCount_T_184 = _zeroCount_T_183 + _GEN_4317; // @[BufferAMSNew.scala 38:70]
  wire [14:0] _GEN_4318 = {{14'd0}, io_adcValues_94 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [15:0] _zeroCount_T_185 = _zeroCount_T_184 + _GEN_4318; // @[BufferAMSNew.scala 38:70]
  wire [15:0] _GEN_4319 = {{15'd0}, io_adcValues_95 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [16:0] zeroCount_5 = _zeroCount_T_185 + _GEN_4319; // @[BufferAMSNew.scala 38:70]
  wire [16:0] _GEN_4320 = {{9'd0}, zeroAccumulators_5}; // @[BufferAMSNew.scala 41:50]
  wire [16:0] _zeroAccumulators_5_T_1 = _GEN_4320 + zeroCount_5; // @[BufferAMSNew.scala 41:50]
  wire [1:0] _zeroCount_T_202 = {{1'd0}, io_adcValues_96 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [1:0] _GEN_4321 = {{1'd0}, io_adcValues_97 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [2:0] _zeroCount_T_203 = _zeroCount_T_202 + _GEN_4321; // @[BufferAMSNew.scala 38:70]
  wire [2:0] _GEN_4322 = {{2'd0}, io_adcValues_98 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [3:0] _zeroCount_T_204 = _zeroCount_T_203 + _GEN_4322; // @[BufferAMSNew.scala 38:70]
  wire [3:0] _GEN_4323 = {{3'd0}, io_adcValues_99 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [4:0] _zeroCount_T_205 = _zeroCount_T_204 + _GEN_4323; // @[BufferAMSNew.scala 38:70]
  wire [4:0] _GEN_4324 = {{4'd0}, io_adcValues_100 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [5:0] _zeroCount_T_206 = _zeroCount_T_205 + _GEN_4324; // @[BufferAMSNew.scala 38:70]
  wire [5:0] _GEN_4325 = {{5'd0}, io_adcValues_101 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [6:0] _zeroCount_T_207 = _zeroCount_T_206 + _GEN_4325; // @[BufferAMSNew.scala 38:70]
  wire [6:0] _GEN_4326 = {{6'd0}, io_adcValues_102 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [7:0] _zeroCount_T_208 = _zeroCount_T_207 + _GEN_4326; // @[BufferAMSNew.scala 38:70]
  wire [7:0] _GEN_4327 = {{7'd0}, io_adcValues_103 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [8:0] _zeroCount_T_209 = _zeroCount_T_208 + _GEN_4327; // @[BufferAMSNew.scala 38:70]
  wire [8:0] _GEN_4328 = {{8'd0}, io_adcValues_104 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [9:0] _zeroCount_T_210 = _zeroCount_T_209 + _GEN_4328; // @[BufferAMSNew.scala 38:70]
  wire [9:0] _GEN_4329 = {{9'd0}, io_adcValues_105 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [10:0] _zeroCount_T_211 = _zeroCount_T_210 + _GEN_4329; // @[BufferAMSNew.scala 38:70]
  wire [10:0] _GEN_4330 = {{10'd0}, io_adcValues_106 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [11:0] _zeroCount_T_212 = _zeroCount_T_211 + _GEN_4330; // @[BufferAMSNew.scala 38:70]
  wire [11:0] _GEN_4331 = {{11'd0}, io_adcValues_107 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [12:0] _zeroCount_T_213 = _zeroCount_T_212 + _GEN_4331; // @[BufferAMSNew.scala 38:70]
  wire [12:0] _GEN_4332 = {{12'd0}, io_adcValues_108 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [13:0] _zeroCount_T_214 = _zeroCount_T_213 + _GEN_4332; // @[BufferAMSNew.scala 38:70]
  wire [13:0] _GEN_4333 = {{13'd0}, io_adcValues_109 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [14:0] _zeroCount_T_215 = _zeroCount_T_214 + _GEN_4333; // @[BufferAMSNew.scala 38:70]
  wire [14:0] _GEN_4334 = {{14'd0}, io_adcValues_110 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [15:0] _zeroCount_T_216 = _zeroCount_T_215 + _GEN_4334; // @[BufferAMSNew.scala 38:70]
  wire [15:0] _GEN_4335 = {{15'd0}, io_adcValues_111 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [16:0] zeroCount_6 = _zeroCount_T_216 + _GEN_4335; // @[BufferAMSNew.scala 38:70]
  wire [16:0] _GEN_4336 = {{9'd0}, zeroAccumulators_6}; // @[BufferAMSNew.scala 41:50]
  wire [16:0] _zeroAccumulators_6_T_1 = _GEN_4336 + zeroCount_6; // @[BufferAMSNew.scala 41:50]
  wire [1:0] _zeroCount_T_233 = {{1'd0}, io_adcValues_112 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [1:0] _GEN_4337 = {{1'd0}, io_adcValues_113 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [2:0] _zeroCount_T_234 = _zeroCount_T_233 + _GEN_4337; // @[BufferAMSNew.scala 38:70]
  wire [2:0] _GEN_4338 = {{2'd0}, io_adcValues_114 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [3:0] _zeroCount_T_235 = _zeroCount_T_234 + _GEN_4338; // @[BufferAMSNew.scala 38:70]
  wire [3:0] _GEN_4339 = {{3'd0}, io_adcValues_115 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [4:0] _zeroCount_T_236 = _zeroCount_T_235 + _GEN_4339; // @[BufferAMSNew.scala 38:70]
  wire [4:0] _GEN_4340 = {{4'd0}, io_adcValues_116 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [5:0] _zeroCount_T_237 = _zeroCount_T_236 + _GEN_4340; // @[BufferAMSNew.scala 38:70]
  wire [5:0] _GEN_4341 = {{5'd0}, io_adcValues_117 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [6:0] _zeroCount_T_238 = _zeroCount_T_237 + _GEN_4341; // @[BufferAMSNew.scala 38:70]
  wire [6:0] _GEN_4342 = {{6'd0}, io_adcValues_118 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [7:0] _zeroCount_T_239 = _zeroCount_T_238 + _GEN_4342; // @[BufferAMSNew.scala 38:70]
  wire [7:0] _GEN_4343 = {{7'd0}, io_adcValues_119 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [8:0] _zeroCount_T_240 = _zeroCount_T_239 + _GEN_4343; // @[BufferAMSNew.scala 38:70]
  wire [8:0] _GEN_4344 = {{8'd0}, io_adcValues_120 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [9:0] _zeroCount_T_241 = _zeroCount_T_240 + _GEN_4344; // @[BufferAMSNew.scala 38:70]
  wire [9:0] _GEN_4345 = {{9'd0}, io_adcValues_121 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [10:0] _zeroCount_T_242 = _zeroCount_T_241 + _GEN_4345; // @[BufferAMSNew.scala 38:70]
  wire [10:0] _GEN_4346 = {{10'd0}, io_adcValues_122 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [11:0] _zeroCount_T_243 = _zeroCount_T_242 + _GEN_4346; // @[BufferAMSNew.scala 38:70]
  wire [11:0] _GEN_4347 = {{11'd0}, io_adcValues_123 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [12:0] _zeroCount_T_244 = _zeroCount_T_243 + _GEN_4347; // @[BufferAMSNew.scala 38:70]
  wire [12:0] _GEN_4348 = {{12'd0}, io_adcValues_124 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [13:0] _zeroCount_T_245 = _zeroCount_T_244 + _GEN_4348; // @[BufferAMSNew.scala 38:70]
  wire [13:0] _GEN_4349 = {{13'd0}, io_adcValues_125 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [14:0] _zeroCount_T_246 = _zeroCount_T_245 + _GEN_4349; // @[BufferAMSNew.scala 38:70]
  wire [14:0] _GEN_4350 = {{14'd0}, io_adcValues_126 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [15:0] _zeroCount_T_247 = _zeroCount_T_246 + _GEN_4350; // @[BufferAMSNew.scala 38:70]
  wire [15:0] _GEN_4351 = {{15'd0}, io_adcValues_127 == 8'h0}; // @[BufferAMSNew.scala 38:70]
  wire [16:0] zeroCount_7 = _zeroCount_T_247 + _GEN_4351; // @[BufferAMSNew.scala 38:70]
  wire [16:0] _GEN_4352 = {{9'd0}, zeroAccumulators_7}; // @[BufferAMSNew.scala 41:50]
  wire [16:0] _zeroAccumulators_7_T_1 = _GEN_4352 + zeroCount_7; // @[BufferAMSNew.scala 41:50]
  wire [16:0] _GEN_2048 = zeroAccumulators_0 < zeroAccumulators_1 ? {{9'd0}, zeroAccumulators_1} :
    _zeroAccumulators_0_T_1; // @[BufferAMSNew.scala 41:27 47:61 50:31]
  wire [16:0] _GEN_2049 = zeroAccumulators_0 < zeroAccumulators_1 ? {{9'd0}, zeroAccumulators_0} :
    _zeroAccumulators_1_T_1; // @[BufferAMSNew.scala 41:27 47:61 51:35]
  wire [3:0] _GEN_2050 = zeroAccumulators_0 < zeroAccumulators_1 ? indexAccumulators_1 : indexAccumulators_0; // @[BufferAMSNew.scala 47:61 55:32 17:34]
  wire [3:0] _GEN_2051 = zeroAccumulators_0 < zeroAccumulators_1 ? indexAccumulators_0 : indexAccumulators_1; // @[BufferAMSNew.scala 17:34 47:61 56:36]
  wire [16:0] _GEN_2052 = zeroAccumulators_1 < zeroAccumulators_2 ? {{9'd0}, zeroAccumulators_2} : _GEN_2049; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2053 = zeroAccumulators_1 < zeroAccumulators_2 ? {{9'd0}, zeroAccumulators_1} :
    _zeroAccumulators_2_T_1; // @[BufferAMSNew.scala 41:27 47:61 51:35]
  wire [3:0] _GEN_2054 = zeroAccumulators_1 < zeroAccumulators_2 ? indexAccumulators_2 : _GEN_2051; // @[BufferAMSNew.scala 47:61 55:32]
  wire [3:0] _GEN_2055 = zeroAccumulators_1 < zeroAccumulators_2 ? indexAccumulators_1 : indexAccumulators_2; // @[BufferAMSNew.scala 17:34 47:61 56:36]
  wire [16:0] _GEN_2056 = zeroAccumulators_2 < zeroAccumulators_3 ? {{9'd0}, zeroAccumulators_3} : _GEN_2053; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2057 = zeroAccumulators_2 < zeroAccumulators_3 ? {{9'd0}, zeroAccumulators_2} :
    _zeroAccumulators_3_T_1; // @[BufferAMSNew.scala 41:27 47:61 51:35]
  wire [3:0] _GEN_2058 = zeroAccumulators_2 < zeroAccumulators_3 ? indexAccumulators_3 : _GEN_2055; // @[BufferAMSNew.scala 47:61 55:32]
  wire [3:0] _GEN_2059 = zeroAccumulators_2 < zeroAccumulators_3 ? indexAccumulators_2 : indexAccumulators_3; // @[BufferAMSNew.scala 17:34 47:61 56:36]
  wire [16:0] _GEN_2060 = zeroAccumulators_3 < zeroAccumulators_4 ? {{9'd0}, zeroAccumulators_4} : _GEN_2057; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2061 = zeroAccumulators_3 < zeroAccumulators_4 ? {{9'd0}, zeroAccumulators_3} :
    _zeroAccumulators_4_T_1; // @[BufferAMSNew.scala 41:27 47:61 51:35]
  wire [3:0] _GEN_2062 = zeroAccumulators_3 < zeroAccumulators_4 ? indexAccumulators_4 : _GEN_2059; // @[BufferAMSNew.scala 47:61 55:32]
  wire [3:0] _GEN_2063 = zeroAccumulators_3 < zeroAccumulators_4 ? indexAccumulators_3 : indexAccumulators_4; // @[BufferAMSNew.scala 17:34 47:61 56:36]
  wire [16:0] _GEN_2064 = zeroAccumulators_4 < zeroAccumulators_5 ? {{9'd0}, zeroAccumulators_5} : _GEN_2061; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2065 = zeroAccumulators_4 < zeroAccumulators_5 ? {{9'd0}, zeroAccumulators_4} :
    _zeroAccumulators_5_T_1; // @[BufferAMSNew.scala 41:27 47:61 51:35]
  wire [3:0] _GEN_2066 = zeroAccumulators_4 < zeroAccumulators_5 ? indexAccumulators_5 : _GEN_2063; // @[BufferAMSNew.scala 47:61 55:32]
  wire [3:0] _GEN_2067 = zeroAccumulators_4 < zeroAccumulators_5 ? indexAccumulators_4 : indexAccumulators_5; // @[BufferAMSNew.scala 17:34 47:61 56:36]
  wire [16:0] _GEN_2068 = zeroAccumulators_5 < zeroAccumulators_6 ? {{9'd0}, zeroAccumulators_6} : _GEN_2065; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2069 = zeroAccumulators_5 < zeroAccumulators_6 ? {{9'd0}, zeroAccumulators_5} :
    _zeroAccumulators_6_T_1; // @[BufferAMSNew.scala 41:27 47:61 51:35]
  wire [3:0] _GEN_2070 = zeroAccumulators_5 < zeroAccumulators_6 ? indexAccumulators_6 : _GEN_2067; // @[BufferAMSNew.scala 47:61 55:32]
  wire [3:0] _GEN_2071 = zeroAccumulators_5 < zeroAccumulators_6 ? indexAccumulators_5 : indexAccumulators_6; // @[BufferAMSNew.scala 17:34 47:61 56:36]
  wire [16:0] _GEN_2072 = zeroAccumulators_6 < zeroAccumulators_7 ? {{9'd0}, zeroAccumulators_7} : _GEN_2069; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2073 = zeroAccumulators_6 < zeroAccumulators_7 ? {{9'd0}, zeroAccumulators_6} :
    _zeroAccumulators_7_T_1; // @[BufferAMSNew.scala 41:27 47:61 51:35]
  wire [16:0] _GEN_2076 = zeroAccumulators_0 < zeroAccumulators_1 ? {{9'd0}, zeroAccumulators_1} : _GEN_2048; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2077 = zeroAccumulators_0 < zeroAccumulators_1 ? {{9'd0}, zeroAccumulators_0} : _GEN_2052; // @[BufferAMSNew.scala 47:61 51:35]
  wire [3:0] _GEN_2078 = zeroAccumulators_0 < zeroAccumulators_1 ? indexAccumulators_1 : _GEN_2050; // @[BufferAMSNew.scala 47:61 55:32]
  wire [3:0] _GEN_2079 = zeroAccumulators_0 < zeroAccumulators_1 ? indexAccumulators_0 : _GEN_2054; // @[BufferAMSNew.scala 47:61 56:36]
  wire [16:0] _GEN_2080 = zeroAccumulators_1 < zeroAccumulators_2 ? {{9'd0}, zeroAccumulators_2} : _GEN_2077; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2081 = zeroAccumulators_1 < zeroAccumulators_2 ? {{9'd0}, zeroAccumulators_1} : _GEN_2056; // @[BufferAMSNew.scala 47:61 51:35]
  wire [3:0] _GEN_2082 = zeroAccumulators_1 < zeroAccumulators_2 ? indexAccumulators_2 : _GEN_2079; // @[BufferAMSNew.scala 47:61 55:32]
  wire [3:0] _GEN_2083 = zeroAccumulators_1 < zeroAccumulators_2 ? indexAccumulators_1 : _GEN_2058; // @[BufferAMSNew.scala 47:61 56:36]
  wire [16:0] _GEN_2084 = zeroAccumulators_2 < zeroAccumulators_3 ? {{9'd0}, zeroAccumulators_3} : _GEN_2081; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2085 = zeroAccumulators_2 < zeroAccumulators_3 ? {{9'd0}, zeroAccumulators_2} : _GEN_2060; // @[BufferAMSNew.scala 47:61 51:35]
  wire [3:0] _GEN_2086 = zeroAccumulators_2 < zeroAccumulators_3 ? indexAccumulators_3 : _GEN_2083; // @[BufferAMSNew.scala 47:61 55:32]
  wire [3:0] _GEN_2087 = zeroAccumulators_2 < zeroAccumulators_3 ? indexAccumulators_2 : _GEN_2062; // @[BufferAMSNew.scala 47:61 56:36]
  wire [16:0] _GEN_2088 = zeroAccumulators_3 < zeroAccumulators_4 ? {{9'd0}, zeroAccumulators_4} : _GEN_2085; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2089 = zeroAccumulators_3 < zeroAccumulators_4 ? {{9'd0}, zeroAccumulators_3} : _GEN_2064; // @[BufferAMSNew.scala 47:61 51:35]
  wire [3:0] _GEN_2090 = zeroAccumulators_3 < zeroAccumulators_4 ? indexAccumulators_4 : _GEN_2087; // @[BufferAMSNew.scala 47:61 55:32]
  wire [3:0] _GEN_2091 = zeroAccumulators_3 < zeroAccumulators_4 ? indexAccumulators_3 : _GEN_2066; // @[BufferAMSNew.scala 47:61 56:36]
  wire [16:0] _GEN_2092 = zeroAccumulators_4 < zeroAccumulators_5 ? {{9'd0}, zeroAccumulators_5} : _GEN_2089; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2093 = zeroAccumulators_4 < zeroAccumulators_5 ? {{9'd0}, zeroAccumulators_4} : _GEN_2068; // @[BufferAMSNew.scala 47:61 51:35]
  wire [3:0] _GEN_2094 = zeroAccumulators_4 < zeroAccumulators_5 ? indexAccumulators_5 : _GEN_2091; // @[BufferAMSNew.scala 47:61 55:32]
  wire [3:0] _GEN_2095 = zeroAccumulators_4 < zeroAccumulators_5 ? indexAccumulators_4 : _GEN_2070; // @[BufferAMSNew.scala 47:61 56:36]
  wire [16:0] _GEN_2096 = zeroAccumulators_5 < zeroAccumulators_6 ? {{9'd0}, zeroAccumulators_6} : _GEN_2093; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2097 = zeroAccumulators_5 < zeroAccumulators_6 ? {{9'd0}, zeroAccumulators_5} : _GEN_2072; // @[BufferAMSNew.scala 47:61 51:35]
  wire [16:0] _GEN_2100 = zeroAccumulators_0 < zeroAccumulators_1 ? {{9'd0}, zeroAccumulators_1} : _GEN_2076; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2101 = zeroAccumulators_0 < zeroAccumulators_1 ? {{9'd0}, zeroAccumulators_0} : _GEN_2080; // @[BufferAMSNew.scala 47:61 51:35]
  wire [3:0] _GEN_2102 = zeroAccumulators_0 < zeroAccumulators_1 ? indexAccumulators_1 : _GEN_2078; // @[BufferAMSNew.scala 47:61 55:32]
  wire [3:0] _GEN_2103 = zeroAccumulators_0 < zeroAccumulators_1 ? indexAccumulators_0 : _GEN_2082; // @[BufferAMSNew.scala 47:61 56:36]
  wire [16:0] _GEN_2104 = zeroAccumulators_1 < zeroAccumulators_2 ? {{9'd0}, zeroAccumulators_2} : _GEN_2101; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2105 = zeroAccumulators_1 < zeroAccumulators_2 ? {{9'd0}, zeroAccumulators_1} : _GEN_2084; // @[BufferAMSNew.scala 47:61 51:35]
  wire [3:0] _GEN_2106 = zeroAccumulators_1 < zeroAccumulators_2 ? indexAccumulators_2 : _GEN_2103; // @[BufferAMSNew.scala 47:61 55:32]
  wire [3:0] _GEN_2107 = zeroAccumulators_1 < zeroAccumulators_2 ? indexAccumulators_1 : _GEN_2086; // @[BufferAMSNew.scala 47:61 56:36]
  wire [16:0] _GEN_2108 = zeroAccumulators_2 < zeroAccumulators_3 ? {{9'd0}, zeroAccumulators_3} : _GEN_2105; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2109 = zeroAccumulators_2 < zeroAccumulators_3 ? {{9'd0}, zeroAccumulators_2} : _GEN_2088; // @[BufferAMSNew.scala 47:61 51:35]
  wire [3:0] _GEN_2110 = zeroAccumulators_2 < zeroAccumulators_3 ? indexAccumulators_3 : _GEN_2107; // @[BufferAMSNew.scala 47:61 55:32]
  wire [3:0] _GEN_2111 = zeroAccumulators_2 < zeroAccumulators_3 ? indexAccumulators_2 : _GEN_2090; // @[BufferAMSNew.scala 47:61 56:36]
  wire [16:0] _GEN_2112 = zeroAccumulators_3 < zeroAccumulators_4 ? {{9'd0}, zeroAccumulators_4} : _GEN_2109; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2113 = zeroAccumulators_3 < zeroAccumulators_4 ? {{9'd0}, zeroAccumulators_3} : _GEN_2092; // @[BufferAMSNew.scala 47:61 51:35]
  wire [3:0] _GEN_2114 = zeroAccumulators_3 < zeroAccumulators_4 ? indexAccumulators_4 : _GEN_2111; // @[BufferAMSNew.scala 47:61 55:32]
  wire [3:0] _GEN_2115 = zeroAccumulators_3 < zeroAccumulators_4 ? indexAccumulators_3 : _GEN_2094; // @[BufferAMSNew.scala 47:61 56:36]
  wire [16:0] _GEN_2116 = zeroAccumulators_4 < zeroAccumulators_5 ? {{9'd0}, zeroAccumulators_5} : _GEN_2113; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2117 = zeroAccumulators_4 < zeroAccumulators_5 ? {{9'd0}, zeroAccumulators_4} : _GEN_2096; // @[BufferAMSNew.scala 47:61 51:35]
  wire [16:0] _GEN_2120 = zeroAccumulators_0 < zeroAccumulators_1 ? {{9'd0}, zeroAccumulators_1} : _GEN_2100; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2121 = zeroAccumulators_0 < zeroAccumulators_1 ? {{9'd0}, zeroAccumulators_0} : _GEN_2104; // @[BufferAMSNew.scala 47:61 51:35]
  wire [3:0] _GEN_2122 = zeroAccumulators_0 < zeroAccumulators_1 ? indexAccumulators_1 : _GEN_2102; // @[BufferAMSNew.scala 47:61 55:32]
  wire [3:0] _GEN_2123 = zeroAccumulators_0 < zeroAccumulators_1 ? indexAccumulators_0 : _GEN_2106; // @[BufferAMSNew.scala 47:61 56:36]
  wire [16:0] _GEN_2124 = zeroAccumulators_1 < zeroAccumulators_2 ? {{9'd0}, zeroAccumulators_2} : _GEN_2121; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2125 = zeroAccumulators_1 < zeroAccumulators_2 ? {{9'd0}, zeroAccumulators_1} : _GEN_2108; // @[BufferAMSNew.scala 47:61 51:35]
  wire [3:0] _GEN_2126 = zeroAccumulators_1 < zeroAccumulators_2 ? indexAccumulators_2 : _GEN_2123; // @[BufferAMSNew.scala 47:61 55:32]
  wire [3:0] _GEN_2127 = zeroAccumulators_1 < zeroAccumulators_2 ? indexAccumulators_1 : _GEN_2110; // @[BufferAMSNew.scala 47:61 56:36]
  wire [16:0] _GEN_2128 = zeroAccumulators_2 < zeroAccumulators_3 ? {{9'd0}, zeroAccumulators_3} : _GEN_2125; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2129 = zeroAccumulators_2 < zeroAccumulators_3 ? {{9'd0}, zeroAccumulators_2} : _GEN_2112; // @[BufferAMSNew.scala 47:61 51:35]
  wire [3:0] _GEN_2130 = zeroAccumulators_2 < zeroAccumulators_3 ? indexAccumulators_3 : _GEN_2127; // @[BufferAMSNew.scala 47:61 55:32]
  wire [3:0] _GEN_2131 = zeroAccumulators_2 < zeroAccumulators_3 ? indexAccumulators_2 : _GEN_2114; // @[BufferAMSNew.scala 47:61 56:36]
  wire [16:0] _GEN_2132 = zeroAccumulators_3 < zeroAccumulators_4 ? {{9'd0}, zeroAccumulators_4} : _GEN_2129; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2133 = zeroAccumulators_3 < zeroAccumulators_4 ? {{9'd0}, zeroAccumulators_3} : _GEN_2116; // @[BufferAMSNew.scala 47:61 51:35]
  wire [16:0] _GEN_2136 = zeroAccumulators_0 < zeroAccumulators_1 ? {{9'd0}, zeroAccumulators_1} : _GEN_2120; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2137 = zeroAccumulators_0 < zeroAccumulators_1 ? {{9'd0}, zeroAccumulators_0} : _GEN_2124; // @[BufferAMSNew.scala 47:61 51:35]
  wire [3:0] _GEN_2138 = zeroAccumulators_0 < zeroAccumulators_1 ? indexAccumulators_1 : _GEN_2122; // @[BufferAMSNew.scala 47:61 55:32]
  wire [3:0] _GEN_2139 = zeroAccumulators_0 < zeroAccumulators_1 ? indexAccumulators_0 : _GEN_2126; // @[BufferAMSNew.scala 47:61 56:36]
  wire [16:0] _GEN_2140 = zeroAccumulators_1 < zeroAccumulators_2 ? {{9'd0}, zeroAccumulators_2} : _GEN_2137; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2141 = zeroAccumulators_1 < zeroAccumulators_2 ? {{9'd0}, zeroAccumulators_1} : _GEN_2128; // @[BufferAMSNew.scala 47:61 51:35]
  wire [3:0] _GEN_2142 = zeroAccumulators_1 < zeroAccumulators_2 ? indexAccumulators_2 : _GEN_2139; // @[BufferAMSNew.scala 47:61 55:32]
  wire [3:0] _GEN_2143 = zeroAccumulators_1 < zeroAccumulators_2 ? indexAccumulators_1 : _GEN_2130; // @[BufferAMSNew.scala 47:61 56:36]
  wire [16:0] _GEN_2144 = zeroAccumulators_2 < zeroAccumulators_3 ? {{9'd0}, zeroAccumulators_3} : _GEN_2141; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2145 = zeroAccumulators_2 < zeroAccumulators_3 ? {{9'd0}, zeroAccumulators_2} : _GEN_2132; // @[BufferAMSNew.scala 47:61 51:35]
  wire [16:0] _GEN_2148 = zeroAccumulators_0 < zeroAccumulators_1 ? {{9'd0}, zeroAccumulators_1} : _GEN_2136; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2149 = zeroAccumulators_0 < zeroAccumulators_1 ? {{9'd0}, zeroAccumulators_0} : _GEN_2140; // @[BufferAMSNew.scala 47:61 51:35]
  wire [3:0] _GEN_2151 = zeroAccumulators_0 < zeroAccumulators_1 ? indexAccumulators_0 : _GEN_2142; // @[BufferAMSNew.scala 47:61 56:36]
  wire [16:0] _GEN_2152 = zeroAccumulators_1 < zeroAccumulators_2 ? {{9'd0}, zeroAccumulators_2} : _GEN_2149; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2153 = zeroAccumulators_1 < zeroAccumulators_2 ? {{9'd0}, zeroAccumulators_1} : _GEN_2144; // @[BufferAMSNew.scala 47:61 51:35]
  wire [16:0] _GEN_2156 = zeroAccumulators_0 < zeroAccumulators_1 ? {{9'd0}, zeroAccumulators_1} : _GEN_2148; // @[BufferAMSNew.scala 47:61 50:31]
  wire [16:0] _GEN_2157 = zeroAccumulators_0 < zeroAccumulators_1 ? {{9'd0}, zeroAccumulators_0} : _GEN_2152; // @[BufferAMSNew.scala 47:61 51:35]
  wire [16:0] _GEN_2161 = lineCounter == 4'hf ? 17'h0 : _GEN_2156; // @[BufferAMSNew.scala 28:30 30:22]
  wire [16:0] _GEN_2162 = lineCounter == 4'hf ? 17'h0 : _GEN_2157; // @[BufferAMSNew.scala 28:30 30:22]
  wire [16:0] _GEN_2163 = lineCounter == 4'hf ? 17'h0 : _GEN_2153; // @[BufferAMSNew.scala 28:30 30:22]
  wire [16:0] _GEN_2164 = lineCounter == 4'hf ? 17'h0 : _GEN_2145; // @[BufferAMSNew.scala 28:30 30:22]
  wire [16:0] _GEN_2165 = lineCounter == 4'hf ? 17'h0 : _GEN_2133; // @[BufferAMSNew.scala 28:30 30:22]
  wire [16:0] _GEN_2166 = lineCounter == 4'hf ? 17'h0 : _GEN_2117; // @[BufferAMSNew.scala 28:30 30:22]
  wire [16:0] _GEN_2167 = lineCounter == 4'hf ? 17'h0 : _GEN_2097; // @[BufferAMSNew.scala 28:30 30:22]
  wire [16:0] _GEN_2168 = lineCounter == 4'hf ? 17'h0 : _GEN_2073; // @[BufferAMSNew.scala 28:30 30:22]
  wire [7:0] _GEN_2178 = 4'h1 == lineCounter ? frameBuffer_1_0 : frameBuffer_0_0; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2179 = 4'h2 == lineCounter ? frameBuffer_2_0 : _GEN_2178; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2180 = 4'h3 == lineCounter ? frameBuffer_3_0 : _GEN_2179; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2181 = 4'h4 == lineCounter ? frameBuffer_4_0 : _GEN_2180; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2182 = 4'h5 == lineCounter ? frameBuffer_5_0 : _GEN_2181; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2183 = 4'h6 == lineCounter ? frameBuffer_6_0 : _GEN_2182; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2184 = 4'h7 == lineCounter ? frameBuffer_7_0 : _GEN_2183; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2185 = 4'h8 == lineCounter ? frameBuffer_8_0 : _GEN_2184; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2186 = 4'h9 == lineCounter ? frameBuffer_9_0 : _GEN_2185; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2187 = 4'ha == lineCounter ? frameBuffer_10_0 : _GEN_2186; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2188 = 4'hb == lineCounter ? frameBuffer_11_0 : _GEN_2187; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2189 = 4'hc == lineCounter ? frameBuffer_12_0 : _GEN_2188; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2190 = 4'hd == lineCounter ? frameBuffer_13_0 : _GEN_2189; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2191 = 4'he == lineCounter ? frameBuffer_14_0 : _GEN_2190; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2194 = 4'h1 == lineCounter ? frameBuffer_1_1 : frameBuffer_0_1; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2195 = 4'h2 == lineCounter ? frameBuffer_2_1 : _GEN_2194; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2196 = 4'h3 == lineCounter ? frameBuffer_3_1 : _GEN_2195; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2197 = 4'h4 == lineCounter ? frameBuffer_4_1 : _GEN_2196; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2198 = 4'h5 == lineCounter ? frameBuffer_5_1 : _GEN_2197; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2199 = 4'h6 == lineCounter ? frameBuffer_6_1 : _GEN_2198; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2200 = 4'h7 == lineCounter ? frameBuffer_7_1 : _GEN_2199; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2201 = 4'h8 == lineCounter ? frameBuffer_8_1 : _GEN_2200; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2202 = 4'h9 == lineCounter ? frameBuffer_9_1 : _GEN_2201; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2203 = 4'ha == lineCounter ? frameBuffer_10_1 : _GEN_2202; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2204 = 4'hb == lineCounter ? frameBuffer_11_1 : _GEN_2203; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2205 = 4'hc == lineCounter ? frameBuffer_12_1 : _GEN_2204; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2206 = 4'hd == lineCounter ? frameBuffer_13_1 : _GEN_2205; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2207 = 4'he == lineCounter ? frameBuffer_14_1 : _GEN_2206; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2210 = 4'h1 == lineCounter ? frameBuffer_1_2 : frameBuffer_0_2; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2211 = 4'h2 == lineCounter ? frameBuffer_2_2 : _GEN_2210; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2212 = 4'h3 == lineCounter ? frameBuffer_3_2 : _GEN_2211; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2213 = 4'h4 == lineCounter ? frameBuffer_4_2 : _GEN_2212; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2214 = 4'h5 == lineCounter ? frameBuffer_5_2 : _GEN_2213; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2215 = 4'h6 == lineCounter ? frameBuffer_6_2 : _GEN_2214; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2216 = 4'h7 == lineCounter ? frameBuffer_7_2 : _GEN_2215; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2217 = 4'h8 == lineCounter ? frameBuffer_8_2 : _GEN_2216; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2218 = 4'h9 == lineCounter ? frameBuffer_9_2 : _GEN_2217; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2219 = 4'ha == lineCounter ? frameBuffer_10_2 : _GEN_2218; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2220 = 4'hb == lineCounter ? frameBuffer_11_2 : _GEN_2219; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2221 = 4'hc == lineCounter ? frameBuffer_12_2 : _GEN_2220; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2222 = 4'hd == lineCounter ? frameBuffer_13_2 : _GEN_2221; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2223 = 4'he == lineCounter ? frameBuffer_14_2 : _GEN_2222; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2226 = 4'h1 == lineCounter ? frameBuffer_1_3 : frameBuffer_0_3; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2227 = 4'h2 == lineCounter ? frameBuffer_2_3 : _GEN_2226; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2228 = 4'h3 == lineCounter ? frameBuffer_3_3 : _GEN_2227; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2229 = 4'h4 == lineCounter ? frameBuffer_4_3 : _GEN_2228; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2230 = 4'h5 == lineCounter ? frameBuffer_5_3 : _GEN_2229; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2231 = 4'h6 == lineCounter ? frameBuffer_6_3 : _GEN_2230; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2232 = 4'h7 == lineCounter ? frameBuffer_7_3 : _GEN_2231; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2233 = 4'h8 == lineCounter ? frameBuffer_8_3 : _GEN_2232; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2234 = 4'h9 == lineCounter ? frameBuffer_9_3 : _GEN_2233; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2235 = 4'ha == lineCounter ? frameBuffer_10_3 : _GEN_2234; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2236 = 4'hb == lineCounter ? frameBuffer_11_3 : _GEN_2235; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2237 = 4'hc == lineCounter ? frameBuffer_12_3 : _GEN_2236; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2238 = 4'hd == lineCounter ? frameBuffer_13_3 : _GEN_2237; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2239 = 4'he == lineCounter ? frameBuffer_14_3 : _GEN_2238; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2242 = 4'h1 == lineCounter ? frameBuffer_1_4 : frameBuffer_0_4; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2243 = 4'h2 == lineCounter ? frameBuffer_2_4 : _GEN_2242; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2244 = 4'h3 == lineCounter ? frameBuffer_3_4 : _GEN_2243; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2245 = 4'h4 == lineCounter ? frameBuffer_4_4 : _GEN_2244; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2246 = 4'h5 == lineCounter ? frameBuffer_5_4 : _GEN_2245; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2247 = 4'h6 == lineCounter ? frameBuffer_6_4 : _GEN_2246; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2248 = 4'h7 == lineCounter ? frameBuffer_7_4 : _GEN_2247; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2249 = 4'h8 == lineCounter ? frameBuffer_8_4 : _GEN_2248; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2250 = 4'h9 == lineCounter ? frameBuffer_9_4 : _GEN_2249; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2251 = 4'ha == lineCounter ? frameBuffer_10_4 : _GEN_2250; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2252 = 4'hb == lineCounter ? frameBuffer_11_4 : _GEN_2251; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2253 = 4'hc == lineCounter ? frameBuffer_12_4 : _GEN_2252; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2254 = 4'hd == lineCounter ? frameBuffer_13_4 : _GEN_2253; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2255 = 4'he == lineCounter ? frameBuffer_14_4 : _GEN_2254; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2258 = 4'h1 == lineCounter ? frameBuffer_1_5 : frameBuffer_0_5; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2259 = 4'h2 == lineCounter ? frameBuffer_2_5 : _GEN_2258; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2260 = 4'h3 == lineCounter ? frameBuffer_3_5 : _GEN_2259; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2261 = 4'h4 == lineCounter ? frameBuffer_4_5 : _GEN_2260; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2262 = 4'h5 == lineCounter ? frameBuffer_5_5 : _GEN_2261; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2263 = 4'h6 == lineCounter ? frameBuffer_6_5 : _GEN_2262; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2264 = 4'h7 == lineCounter ? frameBuffer_7_5 : _GEN_2263; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2265 = 4'h8 == lineCounter ? frameBuffer_8_5 : _GEN_2264; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2266 = 4'h9 == lineCounter ? frameBuffer_9_5 : _GEN_2265; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2267 = 4'ha == lineCounter ? frameBuffer_10_5 : _GEN_2266; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2268 = 4'hb == lineCounter ? frameBuffer_11_5 : _GEN_2267; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2269 = 4'hc == lineCounter ? frameBuffer_12_5 : _GEN_2268; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2270 = 4'hd == lineCounter ? frameBuffer_13_5 : _GEN_2269; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2271 = 4'he == lineCounter ? frameBuffer_14_5 : _GEN_2270; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2274 = 4'h1 == lineCounter ? frameBuffer_1_6 : frameBuffer_0_6; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2275 = 4'h2 == lineCounter ? frameBuffer_2_6 : _GEN_2274; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2276 = 4'h3 == lineCounter ? frameBuffer_3_6 : _GEN_2275; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2277 = 4'h4 == lineCounter ? frameBuffer_4_6 : _GEN_2276; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2278 = 4'h5 == lineCounter ? frameBuffer_5_6 : _GEN_2277; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2279 = 4'h6 == lineCounter ? frameBuffer_6_6 : _GEN_2278; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2280 = 4'h7 == lineCounter ? frameBuffer_7_6 : _GEN_2279; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2281 = 4'h8 == lineCounter ? frameBuffer_8_6 : _GEN_2280; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2282 = 4'h9 == lineCounter ? frameBuffer_9_6 : _GEN_2281; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2283 = 4'ha == lineCounter ? frameBuffer_10_6 : _GEN_2282; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2284 = 4'hb == lineCounter ? frameBuffer_11_6 : _GEN_2283; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2285 = 4'hc == lineCounter ? frameBuffer_12_6 : _GEN_2284; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2286 = 4'hd == lineCounter ? frameBuffer_13_6 : _GEN_2285; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2287 = 4'he == lineCounter ? frameBuffer_14_6 : _GEN_2286; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2290 = 4'h1 == lineCounter ? frameBuffer_1_7 : frameBuffer_0_7; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2291 = 4'h2 == lineCounter ? frameBuffer_2_7 : _GEN_2290; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2292 = 4'h3 == lineCounter ? frameBuffer_3_7 : _GEN_2291; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2293 = 4'h4 == lineCounter ? frameBuffer_4_7 : _GEN_2292; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2294 = 4'h5 == lineCounter ? frameBuffer_5_7 : _GEN_2293; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2295 = 4'h6 == lineCounter ? frameBuffer_6_7 : _GEN_2294; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2296 = 4'h7 == lineCounter ? frameBuffer_7_7 : _GEN_2295; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2297 = 4'h8 == lineCounter ? frameBuffer_8_7 : _GEN_2296; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2298 = 4'h9 == lineCounter ? frameBuffer_9_7 : _GEN_2297; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2299 = 4'ha == lineCounter ? frameBuffer_10_7 : _GEN_2298; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2300 = 4'hb == lineCounter ? frameBuffer_11_7 : _GEN_2299; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2301 = 4'hc == lineCounter ? frameBuffer_12_7 : _GEN_2300; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2302 = 4'hd == lineCounter ? frameBuffer_13_7 : _GEN_2301; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2303 = 4'he == lineCounter ? frameBuffer_14_7 : _GEN_2302; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2306 = 4'h1 == lineCounter ? frameBuffer_1_8 : frameBuffer_0_8; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2307 = 4'h2 == lineCounter ? frameBuffer_2_8 : _GEN_2306; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2308 = 4'h3 == lineCounter ? frameBuffer_3_8 : _GEN_2307; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2309 = 4'h4 == lineCounter ? frameBuffer_4_8 : _GEN_2308; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2310 = 4'h5 == lineCounter ? frameBuffer_5_8 : _GEN_2309; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2311 = 4'h6 == lineCounter ? frameBuffer_6_8 : _GEN_2310; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2312 = 4'h7 == lineCounter ? frameBuffer_7_8 : _GEN_2311; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2313 = 4'h8 == lineCounter ? frameBuffer_8_8 : _GEN_2312; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2314 = 4'h9 == lineCounter ? frameBuffer_9_8 : _GEN_2313; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2315 = 4'ha == lineCounter ? frameBuffer_10_8 : _GEN_2314; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2316 = 4'hb == lineCounter ? frameBuffer_11_8 : _GEN_2315; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2317 = 4'hc == lineCounter ? frameBuffer_12_8 : _GEN_2316; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2318 = 4'hd == lineCounter ? frameBuffer_13_8 : _GEN_2317; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2319 = 4'he == lineCounter ? frameBuffer_14_8 : _GEN_2318; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2322 = 4'h1 == lineCounter ? frameBuffer_1_9 : frameBuffer_0_9; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2323 = 4'h2 == lineCounter ? frameBuffer_2_9 : _GEN_2322; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2324 = 4'h3 == lineCounter ? frameBuffer_3_9 : _GEN_2323; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2325 = 4'h4 == lineCounter ? frameBuffer_4_9 : _GEN_2324; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2326 = 4'h5 == lineCounter ? frameBuffer_5_9 : _GEN_2325; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2327 = 4'h6 == lineCounter ? frameBuffer_6_9 : _GEN_2326; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2328 = 4'h7 == lineCounter ? frameBuffer_7_9 : _GEN_2327; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2329 = 4'h8 == lineCounter ? frameBuffer_8_9 : _GEN_2328; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2330 = 4'h9 == lineCounter ? frameBuffer_9_9 : _GEN_2329; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2331 = 4'ha == lineCounter ? frameBuffer_10_9 : _GEN_2330; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2332 = 4'hb == lineCounter ? frameBuffer_11_9 : _GEN_2331; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2333 = 4'hc == lineCounter ? frameBuffer_12_9 : _GEN_2332; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2334 = 4'hd == lineCounter ? frameBuffer_13_9 : _GEN_2333; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2335 = 4'he == lineCounter ? frameBuffer_14_9 : _GEN_2334; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2338 = 4'h1 == lineCounter ? frameBuffer_1_10 : frameBuffer_0_10; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2339 = 4'h2 == lineCounter ? frameBuffer_2_10 : _GEN_2338; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2340 = 4'h3 == lineCounter ? frameBuffer_3_10 : _GEN_2339; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2341 = 4'h4 == lineCounter ? frameBuffer_4_10 : _GEN_2340; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2342 = 4'h5 == lineCounter ? frameBuffer_5_10 : _GEN_2341; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2343 = 4'h6 == lineCounter ? frameBuffer_6_10 : _GEN_2342; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2344 = 4'h7 == lineCounter ? frameBuffer_7_10 : _GEN_2343; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2345 = 4'h8 == lineCounter ? frameBuffer_8_10 : _GEN_2344; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2346 = 4'h9 == lineCounter ? frameBuffer_9_10 : _GEN_2345; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2347 = 4'ha == lineCounter ? frameBuffer_10_10 : _GEN_2346; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2348 = 4'hb == lineCounter ? frameBuffer_11_10 : _GEN_2347; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2349 = 4'hc == lineCounter ? frameBuffer_12_10 : _GEN_2348; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2350 = 4'hd == lineCounter ? frameBuffer_13_10 : _GEN_2349; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2351 = 4'he == lineCounter ? frameBuffer_14_10 : _GEN_2350; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2354 = 4'h1 == lineCounter ? frameBuffer_1_11 : frameBuffer_0_11; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2355 = 4'h2 == lineCounter ? frameBuffer_2_11 : _GEN_2354; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2356 = 4'h3 == lineCounter ? frameBuffer_3_11 : _GEN_2355; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2357 = 4'h4 == lineCounter ? frameBuffer_4_11 : _GEN_2356; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2358 = 4'h5 == lineCounter ? frameBuffer_5_11 : _GEN_2357; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2359 = 4'h6 == lineCounter ? frameBuffer_6_11 : _GEN_2358; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2360 = 4'h7 == lineCounter ? frameBuffer_7_11 : _GEN_2359; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2361 = 4'h8 == lineCounter ? frameBuffer_8_11 : _GEN_2360; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2362 = 4'h9 == lineCounter ? frameBuffer_9_11 : _GEN_2361; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2363 = 4'ha == lineCounter ? frameBuffer_10_11 : _GEN_2362; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2364 = 4'hb == lineCounter ? frameBuffer_11_11 : _GEN_2363; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2365 = 4'hc == lineCounter ? frameBuffer_12_11 : _GEN_2364; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2366 = 4'hd == lineCounter ? frameBuffer_13_11 : _GEN_2365; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2367 = 4'he == lineCounter ? frameBuffer_14_11 : _GEN_2366; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2370 = 4'h1 == lineCounter ? frameBuffer_1_12 : frameBuffer_0_12; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2371 = 4'h2 == lineCounter ? frameBuffer_2_12 : _GEN_2370; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2372 = 4'h3 == lineCounter ? frameBuffer_3_12 : _GEN_2371; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2373 = 4'h4 == lineCounter ? frameBuffer_4_12 : _GEN_2372; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2374 = 4'h5 == lineCounter ? frameBuffer_5_12 : _GEN_2373; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2375 = 4'h6 == lineCounter ? frameBuffer_6_12 : _GEN_2374; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2376 = 4'h7 == lineCounter ? frameBuffer_7_12 : _GEN_2375; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2377 = 4'h8 == lineCounter ? frameBuffer_8_12 : _GEN_2376; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2378 = 4'h9 == lineCounter ? frameBuffer_9_12 : _GEN_2377; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2379 = 4'ha == lineCounter ? frameBuffer_10_12 : _GEN_2378; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2380 = 4'hb == lineCounter ? frameBuffer_11_12 : _GEN_2379; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2381 = 4'hc == lineCounter ? frameBuffer_12_12 : _GEN_2380; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2382 = 4'hd == lineCounter ? frameBuffer_13_12 : _GEN_2381; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2383 = 4'he == lineCounter ? frameBuffer_14_12 : _GEN_2382; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2386 = 4'h1 == lineCounter ? frameBuffer_1_13 : frameBuffer_0_13; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2387 = 4'h2 == lineCounter ? frameBuffer_2_13 : _GEN_2386; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2388 = 4'h3 == lineCounter ? frameBuffer_3_13 : _GEN_2387; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2389 = 4'h4 == lineCounter ? frameBuffer_4_13 : _GEN_2388; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2390 = 4'h5 == lineCounter ? frameBuffer_5_13 : _GEN_2389; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2391 = 4'h6 == lineCounter ? frameBuffer_6_13 : _GEN_2390; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2392 = 4'h7 == lineCounter ? frameBuffer_7_13 : _GEN_2391; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2393 = 4'h8 == lineCounter ? frameBuffer_8_13 : _GEN_2392; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2394 = 4'h9 == lineCounter ? frameBuffer_9_13 : _GEN_2393; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2395 = 4'ha == lineCounter ? frameBuffer_10_13 : _GEN_2394; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2396 = 4'hb == lineCounter ? frameBuffer_11_13 : _GEN_2395; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2397 = 4'hc == lineCounter ? frameBuffer_12_13 : _GEN_2396; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2398 = 4'hd == lineCounter ? frameBuffer_13_13 : _GEN_2397; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2399 = 4'he == lineCounter ? frameBuffer_14_13 : _GEN_2398; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2402 = 4'h1 == lineCounter ? frameBuffer_1_14 : frameBuffer_0_14; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2403 = 4'h2 == lineCounter ? frameBuffer_2_14 : _GEN_2402; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2404 = 4'h3 == lineCounter ? frameBuffer_3_14 : _GEN_2403; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2405 = 4'h4 == lineCounter ? frameBuffer_4_14 : _GEN_2404; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2406 = 4'h5 == lineCounter ? frameBuffer_5_14 : _GEN_2405; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2407 = 4'h6 == lineCounter ? frameBuffer_6_14 : _GEN_2406; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2408 = 4'h7 == lineCounter ? frameBuffer_7_14 : _GEN_2407; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2409 = 4'h8 == lineCounter ? frameBuffer_8_14 : _GEN_2408; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2410 = 4'h9 == lineCounter ? frameBuffer_9_14 : _GEN_2409; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2411 = 4'ha == lineCounter ? frameBuffer_10_14 : _GEN_2410; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2412 = 4'hb == lineCounter ? frameBuffer_11_14 : _GEN_2411; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2413 = 4'hc == lineCounter ? frameBuffer_12_14 : _GEN_2412; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2414 = 4'hd == lineCounter ? frameBuffer_13_14 : _GEN_2413; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2415 = 4'he == lineCounter ? frameBuffer_14_14 : _GEN_2414; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2418 = 4'h1 == lineCounter ? frameBuffer_1_15 : frameBuffer_0_15; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2419 = 4'h2 == lineCounter ? frameBuffer_2_15 : _GEN_2418; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2420 = 4'h3 == lineCounter ? frameBuffer_3_15 : _GEN_2419; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2421 = 4'h4 == lineCounter ? frameBuffer_4_15 : _GEN_2420; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2422 = 4'h5 == lineCounter ? frameBuffer_5_15 : _GEN_2421; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2423 = 4'h6 == lineCounter ? frameBuffer_6_15 : _GEN_2422; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2424 = 4'h7 == lineCounter ? frameBuffer_7_15 : _GEN_2423; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2425 = 4'h8 == lineCounter ? frameBuffer_8_15 : _GEN_2424; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2426 = 4'h9 == lineCounter ? frameBuffer_9_15 : _GEN_2425; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2427 = 4'ha == lineCounter ? frameBuffer_10_15 : _GEN_2426; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2428 = 4'hb == lineCounter ? frameBuffer_11_15 : _GEN_2427; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2429 = 4'hc == lineCounter ? frameBuffer_12_15 : _GEN_2428; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2430 = 4'hd == lineCounter ? frameBuffer_13_15 : _GEN_2429; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2431 = 4'he == lineCounter ? frameBuffer_14_15 : _GEN_2430; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2434 = 4'h1 == lineCounter ? frameBuffer_1_16 : frameBuffer_0_16; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2435 = 4'h2 == lineCounter ? frameBuffer_2_16 : _GEN_2434; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2436 = 4'h3 == lineCounter ? frameBuffer_3_16 : _GEN_2435; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2437 = 4'h4 == lineCounter ? frameBuffer_4_16 : _GEN_2436; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2438 = 4'h5 == lineCounter ? frameBuffer_5_16 : _GEN_2437; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2439 = 4'h6 == lineCounter ? frameBuffer_6_16 : _GEN_2438; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2440 = 4'h7 == lineCounter ? frameBuffer_7_16 : _GEN_2439; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2441 = 4'h8 == lineCounter ? frameBuffer_8_16 : _GEN_2440; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2442 = 4'h9 == lineCounter ? frameBuffer_9_16 : _GEN_2441; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2443 = 4'ha == lineCounter ? frameBuffer_10_16 : _GEN_2442; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2444 = 4'hb == lineCounter ? frameBuffer_11_16 : _GEN_2443; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2445 = 4'hc == lineCounter ? frameBuffer_12_16 : _GEN_2444; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2446 = 4'hd == lineCounter ? frameBuffer_13_16 : _GEN_2445; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2447 = 4'he == lineCounter ? frameBuffer_14_16 : _GEN_2446; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2450 = 4'h1 == lineCounter ? frameBuffer_1_17 : frameBuffer_0_17; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2451 = 4'h2 == lineCounter ? frameBuffer_2_17 : _GEN_2450; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2452 = 4'h3 == lineCounter ? frameBuffer_3_17 : _GEN_2451; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2453 = 4'h4 == lineCounter ? frameBuffer_4_17 : _GEN_2452; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2454 = 4'h5 == lineCounter ? frameBuffer_5_17 : _GEN_2453; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2455 = 4'h6 == lineCounter ? frameBuffer_6_17 : _GEN_2454; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2456 = 4'h7 == lineCounter ? frameBuffer_7_17 : _GEN_2455; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2457 = 4'h8 == lineCounter ? frameBuffer_8_17 : _GEN_2456; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2458 = 4'h9 == lineCounter ? frameBuffer_9_17 : _GEN_2457; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2459 = 4'ha == lineCounter ? frameBuffer_10_17 : _GEN_2458; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2460 = 4'hb == lineCounter ? frameBuffer_11_17 : _GEN_2459; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2461 = 4'hc == lineCounter ? frameBuffer_12_17 : _GEN_2460; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2462 = 4'hd == lineCounter ? frameBuffer_13_17 : _GEN_2461; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2463 = 4'he == lineCounter ? frameBuffer_14_17 : _GEN_2462; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2466 = 4'h1 == lineCounter ? frameBuffer_1_18 : frameBuffer_0_18; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2467 = 4'h2 == lineCounter ? frameBuffer_2_18 : _GEN_2466; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2468 = 4'h3 == lineCounter ? frameBuffer_3_18 : _GEN_2467; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2469 = 4'h4 == lineCounter ? frameBuffer_4_18 : _GEN_2468; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2470 = 4'h5 == lineCounter ? frameBuffer_5_18 : _GEN_2469; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2471 = 4'h6 == lineCounter ? frameBuffer_6_18 : _GEN_2470; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2472 = 4'h7 == lineCounter ? frameBuffer_7_18 : _GEN_2471; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2473 = 4'h8 == lineCounter ? frameBuffer_8_18 : _GEN_2472; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2474 = 4'h9 == lineCounter ? frameBuffer_9_18 : _GEN_2473; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2475 = 4'ha == lineCounter ? frameBuffer_10_18 : _GEN_2474; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2476 = 4'hb == lineCounter ? frameBuffer_11_18 : _GEN_2475; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2477 = 4'hc == lineCounter ? frameBuffer_12_18 : _GEN_2476; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2478 = 4'hd == lineCounter ? frameBuffer_13_18 : _GEN_2477; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2479 = 4'he == lineCounter ? frameBuffer_14_18 : _GEN_2478; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2482 = 4'h1 == lineCounter ? frameBuffer_1_19 : frameBuffer_0_19; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2483 = 4'h2 == lineCounter ? frameBuffer_2_19 : _GEN_2482; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2484 = 4'h3 == lineCounter ? frameBuffer_3_19 : _GEN_2483; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2485 = 4'h4 == lineCounter ? frameBuffer_4_19 : _GEN_2484; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2486 = 4'h5 == lineCounter ? frameBuffer_5_19 : _GEN_2485; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2487 = 4'h6 == lineCounter ? frameBuffer_6_19 : _GEN_2486; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2488 = 4'h7 == lineCounter ? frameBuffer_7_19 : _GEN_2487; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2489 = 4'h8 == lineCounter ? frameBuffer_8_19 : _GEN_2488; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2490 = 4'h9 == lineCounter ? frameBuffer_9_19 : _GEN_2489; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2491 = 4'ha == lineCounter ? frameBuffer_10_19 : _GEN_2490; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2492 = 4'hb == lineCounter ? frameBuffer_11_19 : _GEN_2491; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2493 = 4'hc == lineCounter ? frameBuffer_12_19 : _GEN_2492; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2494 = 4'hd == lineCounter ? frameBuffer_13_19 : _GEN_2493; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2495 = 4'he == lineCounter ? frameBuffer_14_19 : _GEN_2494; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2498 = 4'h1 == lineCounter ? frameBuffer_1_20 : frameBuffer_0_20; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2499 = 4'h2 == lineCounter ? frameBuffer_2_20 : _GEN_2498; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2500 = 4'h3 == lineCounter ? frameBuffer_3_20 : _GEN_2499; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2501 = 4'h4 == lineCounter ? frameBuffer_4_20 : _GEN_2500; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2502 = 4'h5 == lineCounter ? frameBuffer_5_20 : _GEN_2501; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2503 = 4'h6 == lineCounter ? frameBuffer_6_20 : _GEN_2502; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2504 = 4'h7 == lineCounter ? frameBuffer_7_20 : _GEN_2503; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2505 = 4'h8 == lineCounter ? frameBuffer_8_20 : _GEN_2504; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2506 = 4'h9 == lineCounter ? frameBuffer_9_20 : _GEN_2505; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2507 = 4'ha == lineCounter ? frameBuffer_10_20 : _GEN_2506; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2508 = 4'hb == lineCounter ? frameBuffer_11_20 : _GEN_2507; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2509 = 4'hc == lineCounter ? frameBuffer_12_20 : _GEN_2508; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2510 = 4'hd == lineCounter ? frameBuffer_13_20 : _GEN_2509; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2511 = 4'he == lineCounter ? frameBuffer_14_20 : _GEN_2510; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2514 = 4'h1 == lineCounter ? frameBuffer_1_21 : frameBuffer_0_21; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2515 = 4'h2 == lineCounter ? frameBuffer_2_21 : _GEN_2514; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2516 = 4'h3 == lineCounter ? frameBuffer_3_21 : _GEN_2515; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2517 = 4'h4 == lineCounter ? frameBuffer_4_21 : _GEN_2516; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2518 = 4'h5 == lineCounter ? frameBuffer_5_21 : _GEN_2517; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2519 = 4'h6 == lineCounter ? frameBuffer_6_21 : _GEN_2518; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2520 = 4'h7 == lineCounter ? frameBuffer_7_21 : _GEN_2519; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2521 = 4'h8 == lineCounter ? frameBuffer_8_21 : _GEN_2520; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2522 = 4'h9 == lineCounter ? frameBuffer_9_21 : _GEN_2521; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2523 = 4'ha == lineCounter ? frameBuffer_10_21 : _GEN_2522; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2524 = 4'hb == lineCounter ? frameBuffer_11_21 : _GEN_2523; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2525 = 4'hc == lineCounter ? frameBuffer_12_21 : _GEN_2524; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2526 = 4'hd == lineCounter ? frameBuffer_13_21 : _GEN_2525; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2527 = 4'he == lineCounter ? frameBuffer_14_21 : _GEN_2526; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2530 = 4'h1 == lineCounter ? frameBuffer_1_22 : frameBuffer_0_22; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2531 = 4'h2 == lineCounter ? frameBuffer_2_22 : _GEN_2530; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2532 = 4'h3 == lineCounter ? frameBuffer_3_22 : _GEN_2531; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2533 = 4'h4 == lineCounter ? frameBuffer_4_22 : _GEN_2532; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2534 = 4'h5 == lineCounter ? frameBuffer_5_22 : _GEN_2533; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2535 = 4'h6 == lineCounter ? frameBuffer_6_22 : _GEN_2534; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2536 = 4'h7 == lineCounter ? frameBuffer_7_22 : _GEN_2535; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2537 = 4'h8 == lineCounter ? frameBuffer_8_22 : _GEN_2536; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2538 = 4'h9 == lineCounter ? frameBuffer_9_22 : _GEN_2537; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2539 = 4'ha == lineCounter ? frameBuffer_10_22 : _GEN_2538; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2540 = 4'hb == lineCounter ? frameBuffer_11_22 : _GEN_2539; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2541 = 4'hc == lineCounter ? frameBuffer_12_22 : _GEN_2540; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2542 = 4'hd == lineCounter ? frameBuffer_13_22 : _GEN_2541; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2543 = 4'he == lineCounter ? frameBuffer_14_22 : _GEN_2542; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2546 = 4'h1 == lineCounter ? frameBuffer_1_23 : frameBuffer_0_23; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2547 = 4'h2 == lineCounter ? frameBuffer_2_23 : _GEN_2546; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2548 = 4'h3 == lineCounter ? frameBuffer_3_23 : _GEN_2547; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2549 = 4'h4 == lineCounter ? frameBuffer_4_23 : _GEN_2548; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2550 = 4'h5 == lineCounter ? frameBuffer_5_23 : _GEN_2549; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2551 = 4'h6 == lineCounter ? frameBuffer_6_23 : _GEN_2550; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2552 = 4'h7 == lineCounter ? frameBuffer_7_23 : _GEN_2551; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2553 = 4'h8 == lineCounter ? frameBuffer_8_23 : _GEN_2552; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2554 = 4'h9 == lineCounter ? frameBuffer_9_23 : _GEN_2553; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2555 = 4'ha == lineCounter ? frameBuffer_10_23 : _GEN_2554; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2556 = 4'hb == lineCounter ? frameBuffer_11_23 : _GEN_2555; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2557 = 4'hc == lineCounter ? frameBuffer_12_23 : _GEN_2556; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2558 = 4'hd == lineCounter ? frameBuffer_13_23 : _GEN_2557; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2559 = 4'he == lineCounter ? frameBuffer_14_23 : _GEN_2558; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2562 = 4'h1 == lineCounter ? frameBuffer_1_24 : frameBuffer_0_24; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2563 = 4'h2 == lineCounter ? frameBuffer_2_24 : _GEN_2562; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2564 = 4'h3 == lineCounter ? frameBuffer_3_24 : _GEN_2563; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2565 = 4'h4 == lineCounter ? frameBuffer_4_24 : _GEN_2564; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2566 = 4'h5 == lineCounter ? frameBuffer_5_24 : _GEN_2565; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2567 = 4'h6 == lineCounter ? frameBuffer_6_24 : _GEN_2566; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2568 = 4'h7 == lineCounter ? frameBuffer_7_24 : _GEN_2567; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2569 = 4'h8 == lineCounter ? frameBuffer_8_24 : _GEN_2568; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2570 = 4'h9 == lineCounter ? frameBuffer_9_24 : _GEN_2569; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2571 = 4'ha == lineCounter ? frameBuffer_10_24 : _GEN_2570; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2572 = 4'hb == lineCounter ? frameBuffer_11_24 : _GEN_2571; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2573 = 4'hc == lineCounter ? frameBuffer_12_24 : _GEN_2572; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2574 = 4'hd == lineCounter ? frameBuffer_13_24 : _GEN_2573; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2575 = 4'he == lineCounter ? frameBuffer_14_24 : _GEN_2574; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2578 = 4'h1 == lineCounter ? frameBuffer_1_25 : frameBuffer_0_25; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2579 = 4'h2 == lineCounter ? frameBuffer_2_25 : _GEN_2578; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2580 = 4'h3 == lineCounter ? frameBuffer_3_25 : _GEN_2579; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2581 = 4'h4 == lineCounter ? frameBuffer_4_25 : _GEN_2580; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2582 = 4'h5 == lineCounter ? frameBuffer_5_25 : _GEN_2581; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2583 = 4'h6 == lineCounter ? frameBuffer_6_25 : _GEN_2582; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2584 = 4'h7 == lineCounter ? frameBuffer_7_25 : _GEN_2583; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2585 = 4'h8 == lineCounter ? frameBuffer_8_25 : _GEN_2584; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2586 = 4'h9 == lineCounter ? frameBuffer_9_25 : _GEN_2585; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2587 = 4'ha == lineCounter ? frameBuffer_10_25 : _GEN_2586; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2588 = 4'hb == lineCounter ? frameBuffer_11_25 : _GEN_2587; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2589 = 4'hc == lineCounter ? frameBuffer_12_25 : _GEN_2588; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2590 = 4'hd == lineCounter ? frameBuffer_13_25 : _GEN_2589; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2591 = 4'he == lineCounter ? frameBuffer_14_25 : _GEN_2590; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2594 = 4'h1 == lineCounter ? frameBuffer_1_26 : frameBuffer_0_26; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2595 = 4'h2 == lineCounter ? frameBuffer_2_26 : _GEN_2594; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2596 = 4'h3 == lineCounter ? frameBuffer_3_26 : _GEN_2595; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2597 = 4'h4 == lineCounter ? frameBuffer_4_26 : _GEN_2596; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2598 = 4'h5 == lineCounter ? frameBuffer_5_26 : _GEN_2597; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2599 = 4'h6 == lineCounter ? frameBuffer_6_26 : _GEN_2598; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2600 = 4'h7 == lineCounter ? frameBuffer_7_26 : _GEN_2599; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2601 = 4'h8 == lineCounter ? frameBuffer_8_26 : _GEN_2600; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2602 = 4'h9 == lineCounter ? frameBuffer_9_26 : _GEN_2601; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2603 = 4'ha == lineCounter ? frameBuffer_10_26 : _GEN_2602; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2604 = 4'hb == lineCounter ? frameBuffer_11_26 : _GEN_2603; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2605 = 4'hc == lineCounter ? frameBuffer_12_26 : _GEN_2604; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2606 = 4'hd == lineCounter ? frameBuffer_13_26 : _GEN_2605; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2607 = 4'he == lineCounter ? frameBuffer_14_26 : _GEN_2606; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2610 = 4'h1 == lineCounter ? frameBuffer_1_27 : frameBuffer_0_27; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2611 = 4'h2 == lineCounter ? frameBuffer_2_27 : _GEN_2610; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2612 = 4'h3 == lineCounter ? frameBuffer_3_27 : _GEN_2611; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2613 = 4'h4 == lineCounter ? frameBuffer_4_27 : _GEN_2612; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2614 = 4'h5 == lineCounter ? frameBuffer_5_27 : _GEN_2613; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2615 = 4'h6 == lineCounter ? frameBuffer_6_27 : _GEN_2614; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2616 = 4'h7 == lineCounter ? frameBuffer_7_27 : _GEN_2615; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2617 = 4'h8 == lineCounter ? frameBuffer_8_27 : _GEN_2616; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2618 = 4'h9 == lineCounter ? frameBuffer_9_27 : _GEN_2617; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2619 = 4'ha == lineCounter ? frameBuffer_10_27 : _GEN_2618; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2620 = 4'hb == lineCounter ? frameBuffer_11_27 : _GEN_2619; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2621 = 4'hc == lineCounter ? frameBuffer_12_27 : _GEN_2620; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2622 = 4'hd == lineCounter ? frameBuffer_13_27 : _GEN_2621; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2623 = 4'he == lineCounter ? frameBuffer_14_27 : _GEN_2622; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2626 = 4'h1 == lineCounter ? frameBuffer_1_28 : frameBuffer_0_28; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2627 = 4'h2 == lineCounter ? frameBuffer_2_28 : _GEN_2626; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2628 = 4'h3 == lineCounter ? frameBuffer_3_28 : _GEN_2627; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2629 = 4'h4 == lineCounter ? frameBuffer_4_28 : _GEN_2628; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2630 = 4'h5 == lineCounter ? frameBuffer_5_28 : _GEN_2629; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2631 = 4'h6 == lineCounter ? frameBuffer_6_28 : _GEN_2630; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2632 = 4'h7 == lineCounter ? frameBuffer_7_28 : _GEN_2631; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2633 = 4'h8 == lineCounter ? frameBuffer_8_28 : _GEN_2632; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2634 = 4'h9 == lineCounter ? frameBuffer_9_28 : _GEN_2633; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2635 = 4'ha == lineCounter ? frameBuffer_10_28 : _GEN_2634; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2636 = 4'hb == lineCounter ? frameBuffer_11_28 : _GEN_2635; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2637 = 4'hc == lineCounter ? frameBuffer_12_28 : _GEN_2636; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2638 = 4'hd == lineCounter ? frameBuffer_13_28 : _GEN_2637; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2639 = 4'he == lineCounter ? frameBuffer_14_28 : _GEN_2638; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2642 = 4'h1 == lineCounter ? frameBuffer_1_29 : frameBuffer_0_29; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2643 = 4'h2 == lineCounter ? frameBuffer_2_29 : _GEN_2642; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2644 = 4'h3 == lineCounter ? frameBuffer_3_29 : _GEN_2643; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2645 = 4'h4 == lineCounter ? frameBuffer_4_29 : _GEN_2644; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2646 = 4'h5 == lineCounter ? frameBuffer_5_29 : _GEN_2645; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2647 = 4'h6 == lineCounter ? frameBuffer_6_29 : _GEN_2646; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2648 = 4'h7 == lineCounter ? frameBuffer_7_29 : _GEN_2647; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2649 = 4'h8 == lineCounter ? frameBuffer_8_29 : _GEN_2648; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2650 = 4'h9 == lineCounter ? frameBuffer_9_29 : _GEN_2649; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2651 = 4'ha == lineCounter ? frameBuffer_10_29 : _GEN_2650; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2652 = 4'hb == lineCounter ? frameBuffer_11_29 : _GEN_2651; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2653 = 4'hc == lineCounter ? frameBuffer_12_29 : _GEN_2652; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2654 = 4'hd == lineCounter ? frameBuffer_13_29 : _GEN_2653; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2655 = 4'he == lineCounter ? frameBuffer_14_29 : _GEN_2654; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2658 = 4'h1 == lineCounter ? frameBuffer_1_30 : frameBuffer_0_30; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2659 = 4'h2 == lineCounter ? frameBuffer_2_30 : _GEN_2658; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2660 = 4'h3 == lineCounter ? frameBuffer_3_30 : _GEN_2659; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2661 = 4'h4 == lineCounter ? frameBuffer_4_30 : _GEN_2660; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2662 = 4'h5 == lineCounter ? frameBuffer_5_30 : _GEN_2661; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2663 = 4'h6 == lineCounter ? frameBuffer_6_30 : _GEN_2662; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2664 = 4'h7 == lineCounter ? frameBuffer_7_30 : _GEN_2663; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2665 = 4'h8 == lineCounter ? frameBuffer_8_30 : _GEN_2664; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2666 = 4'h9 == lineCounter ? frameBuffer_9_30 : _GEN_2665; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2667 = 4'ha == lineCounter ? frameBuffer_10_30 : _GEN_2666; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2668 = 4'hb == lineCounter ? frameBuffer_11_30 : _GEN_2667; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2669 = 4'hc == lineCounter ? frameBuffer_12_30 : _GEN_2668; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2670 = 4'hd == lineCounter ? frameBuffer_13_30 : _GEN_2669; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2671 = 4'he == lineCounter ? frameBuffer_14_30 : _GEN_2670; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2674 = 4'h1 == lineCounter ? frameBuffer_1_31 : frameBuffer_0_31; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2675 = 4'h2 == lineCounter ? frameBuffer_2_31 : _GEN_2674; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2676 = 4'h3 == lineCounter ? frameBuffer_3_31 : _GEN_2675; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2677 = 4'h4 == lineCounter ? frameBuffer_4_31 : _GEN_2676; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2678 = 4'h5 == lineCounter ? frameBuffer_5_31 : _GEN_2677; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2679 = 4'h6 == lineCounter ? frameBuffer_6_31 : _GEN_2678; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2680 = 4'h7 == lineCounter ? frameBuffer_7_31 : _GEN_2679; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2681 = 4'h8 == lineCounter ? frameBuffer_8_31 : _GEN_2680; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2682 = 4'h9 == lineCounter ? frameBuffer_9_31 : _GEN_2681; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2683 = 4'ha == lineCounter ? frameBuffer_10_31 : _GEN_2682; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2684 = 4'hb == lineCounter ? frameBuffer_11_31 : _GEN_2683; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2685 = 4'hc == lineCounter ? frameBuffer_12_31 : _GEN_2684; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2686 = 4'hd == lineCounter ? frameBuffer_13_31 : _GEN_2685; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2687 = 4'he == lineCounter ? frameBuffer_14_31 : _GEN_2686; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2690 = 4'h1 == lineCounter ? frameBuffer_1_32 : frameBuffer_0_32; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2691 = 4'h2 == lineCounter ? frameBuffer_2_32 : _GEN_2690; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2692 = 4'h3 == lineCounter ? frameBuffer_3_32 : _GEN_2691; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2693 = 4'h4 == lineCounter ? frameBuffer_4_32 : _GEN_2692; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2694 = 4'h5 == lineCounter ? frameBuffer_5_32 : _GEN_2693; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2695 = 4'h6 == lineCounter ? frameBuffer_6_32 : _GEN_2694; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2696 = 4'h7 == lineCounter ? frameBuffer_7_32 : _GEN_2695; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2697 = 4'h8 == lineCounter ? frameBuffer_8_32 : _GEN_2696; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2698 = 4'h9 == lineCounter ? frameBuffer_9_32 : _GEN_2697; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2699 = 4'ha == lineCounter ? frameBuffer_10_32 : _GEN_2698; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2700 = 4'hb == lineCounter ? frameBuffer_11_32 : _GEN_2699; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2701 = 4'hc == lineCounter ? frameBuffer_12_32 : _GEN_2700; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2702 = 4'hd == lineCounter ? frameBuffer_13_32 : _GEN_2701; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2703 = 4'he == lineCounter ? frameBuffer_14_32 : _GEN_2702; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2706 = 4'h1 == lineCounter ? frameBuffer_1_33 : frameBuffer_0_33; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2707 = 4'h2 == lineCounter ? frameBuffer_2_33 : _GEN_2706; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2708 = 4'h3 == lineCounter ? frameBuffer_3_33 : _GEN_2707; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2709 = 4'h4 == lineCounter ? frameBuffer_4_33 : _GEN_2708; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2710 = 4'h5 == lineCounter ? frameBuffer_5_33 : _GEN_2709; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2711 = 4'h6 == lineCounter ? frameBuffer_6_33 : _GEN_2710; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2712 = 4'h7 == lineCounter ? frameBuffer_7_33 : _GEN_2711; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2713 = 4'h8 == lineCounter ? frameBuffer_8_33 : _GEN_2712; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2714 = 4'h9 == lineCounter ? frameBuffer_9_33 : _GEN_2713; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2715 = 4'ha == lineCounter ? frameBuffer_10_33 : _GEN_2714; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2716 = 4'hb == lineCounter ? frameBuffer_11_33 : _GEN_2715; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2717 = 4'hc == lineCounter ? frameBuffer_12_33 : _GEN_2716; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2718 = 4'hd == lineCounter ? frameBuffer_13_33 : _GEN_2717; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2719 = 4'he == lineCounter ? frameBuffer_14_33 : _GEN_2718; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2722 = 4'h1 == lineCounter ? frameBuffer_1_34 : frameBuffer_0_34; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2723 = 4'h2 == lineCounter ? frameBuffer_2_34 : _GEN_2722; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2724 = 4'h3 == lineCounter ? frameBuffer_3_34 : _GEN_2723; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2725 = 4'h4 == lineCounter ? frameBuffer_4_34 : _GEN_2724; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2726 = 4'h5 == lineCounter ? frameBuffer_5_34 : _GEN_2725; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2727 = 4'h6 == lineCounter ? frameBuffer_6_34 : _GEN_2726; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2728 = 4'h7 == lineCounter ? frameBuffer_7_34 : _GEN_2727; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2729 = 4'h8 == lineCounter ? frameBuffer_8_34 : _GEN_2728; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2730 = 4'h9 == lineCounter ? frameBuffer_9_34 : _GEN_2729; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2731 = 4'ha == lineCounter ? frameBuffer_10_34 : _GEN_2730; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2732 = 4'hb == lineCounter ? frameBuffer_11_34 : _GEN_2731; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2733 = 4'hc == lineCounter ? frameBuffer_12_34 : _GEN_2732; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2734 = 4'hd == lineCounter ? frameBuffer_13_34 : _GEN_2733; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2735 = 4'he == lineCounter ? frameBuffer_14_34 : _GEN_2734; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2738 = 4'h1 == lineCounter ? frameBuffer_1_35 : frameBuffer_0_35; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2739 = 4'h2 == lineCounter ? frameBuffer_2_35 : _GEN_2738; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2740 = 4'h3 == lineCounter ? frameBuffer_3_35 : _GEN_2739; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2741 = 4'h4 == lineCounter ? frameBuffer_4_35 : _GEN_2740; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2742 = 4'h5 == lineCounter ? frameBuffer_5_35 : _GEN_2741; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2743 = 4'h6 == lineCounter ? frameBuffer_6_35 : _GEN_2742; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2744 = 4'h7 == lineCounter ? frameBuffer_7_35 : _GEN_2743; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2745 = 4'h8 == lineCounter ? frameBuffer_8_35 : _GEN_2744; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2746 = 4'h9 == lineCounter ? frameBuffer_9_35 : _GEN_2745; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2747 = 4'ha == lineCounter ? frameBuffer_10_35 : _GEN_2746; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2748 = 4'hb == lineCounter ? frameBuffer_11_35 : _GEN_2747; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2749 = 4'hc == lineCounter ? frameBuffer_12_35 : _GEN_2748; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2750 = 4'hd == lineCounter ? frameBuffer_13_35 : _GEN_2749; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2751 = 4'he == lineCounter ? frameBuffer_14_35 : _GEN_2750; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2754 = 4'h1 == lineCounter ? frameBuffer_1_36 : frameBuffer_0_36; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2755 = 4'h2 == lineCounter ? frameBuffer_2_36 : _GEN_2754; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2756 = 4'h3 == lineCounter ? frameBuffer_3_36 : _GEN_2755; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2757 = 4'h4 == lineCounter ? frameBuffer_4_36 : _GEN_2756; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2758 = 4'h5 == lineCounter ? frameBuffer_5_36 : _GEN_2757; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2759 = 4'h6 == lineCounter ? frameBuffer_6_36 : _GEN_2758; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2760 = 4'h7 == lineCounter ? frameBuffer_7_36 : _GEN_2759; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2761 = 4'h8 == lineCounter ? frameBuffer_8_36 : _GEN_2760; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2762 = 4'h9 == lineCounter ? frameBuffer_9_36 : _GEN_2761; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2763 = 4'ha == lineCounter ? frameBuffer_10_36 : _GEN_2762; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2764 = 4'hb == lineCounter ? frameBuffer_11_36 : _GEN_2763; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2765 = 4'hc == lineCounter ? frameBuffer_12_36 : _GEN_2764; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2766 = 4'hd == lineCounter ? frameBuffer_13_36 : _GEN_2765; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2767 = 4'he == lineCounter ? frameBuffer_14_36 : _GEN_2766; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2770 = 4'h1 == lineCounter ? frameBuffer_1_37 : frameBuffer_0_37; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2771 = 4'h2 == lineCounter ? frameBuffer_2_37 : _GEN_2770; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2772 = 4'h3 == lineCounter ? frameBuffer_3_37 : _GEN_2771; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2773 = 4'h4 == lineCounter ? frameBuffer_4_37 : _GEN_2772; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2774 = 4'h5 == lineCounter ? frameBuffer_5_37 : _GEN_2773; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2775 = 4'h6 == lineCounter ? frameBuffer_6_37 : _GEN_2774; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2776 = 4'h7 == lineCounter ? frameBuffer_7_37 : _GEN_2775; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2777 = 4'h8 == lineCounter ? frameBuffer_8_37 : _GEN_2776; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2778 = 4'h9 == lineCounter ? frameBuffer_9_37 : _GEN_2777; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2779 = 4'ha == lineCounter ? frameBuffer_10_37 : _GEN_2778; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2780 = 4'hb == lineCounter ? frameBuffer_11_37 : _GEN_2779; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2781 = 4'hc == lineCounter ? frameBuffer_12_37 : _GEN_2780; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2782 = 4'hd == lineCounter ? frameBuffer_13_37 : _GEN_2781; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2783 = 4'he == lineCounter ? frameBuffer_14_37 : _GEN_2782; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2786 = 4'h1 == lineCounter ? frameBuffer_1_38 : frameBuffer_0_38; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2787 = 4'h2 == lineCounter ? frameBuffer_2_38 : _GEN_2786; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2788 = 4'h3 == lineCounter ? frameBuffer_3_38 : _GEN_2787; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2789 = 4'h4 == lineCounter ? frameBuffer_4_38 : _GEN_2788; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2790 = 4'h5 == lineCounter ? frameBuffer_5_38 : _GEN_2789; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2791 = 4'h6 == lineCounter ? frameBuffer_6_38 : _GEN_2790; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2792 = 4'h7 == lineCounter ? frameBuffer_7_38 : _GEN_2791; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2793 = 4'h8 == lineCounter ? frameBuffer_8_38 : _GEN_2792; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2794 = 4'h9 == lineCounter ? frameBuffer_9_38 : _GEN_2793; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2795 = 4'ha == lineCounter ? frameBuffer_10_38 : _GEN_2794; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2796 = 4'hb == lineCounter ? frameBuffer_11_38 : _GEN_2795; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2797 = 4'hc == lineCounter ? frameBuffer_12_38 : _GEN_2796; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2798 = 4'hd == lineCounter ? frameBuffer_13_38 : _GEN_2797; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2799 = 4'he == lineCounter ? frameBuffer_14_38 : _GEN_2798; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2802 = 4'h1 == lineCounter ? frameBuffer_1_39 : frameBuffer_0_39; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2803 = 4'h2 == lineCounter ? frameBuffer_2_39 : _GEN_2802; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2804 = 4'h3 == lineCounter ? frameBuffer_3_39 : _GEN_2803; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2805 = 4'h4 == lineCounter ? frameBuffer_4_39 : _GEN_2804; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2806 = 4'h5 == lineCounter ? frameBuffer_5_39 : _GEN_2805; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2807 = 4'h6 == lineCounter ? frameBuffer_6_39 : _GEN_2806; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2808 = 4'h7 == lineCounter ? frameBuffer_7_39 : _GEN_2807; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2809 = 4'h8 == lineCounter ? frameBuffer_8_39 : _GEN_2808; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2810 = 4'h9 == lineCounter ? frameBuffer_9_39 : _GEN_2809; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2811 = 4'ha == lineCounter ? frameBuffer_10_39 : _GEN_2810; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2812 = 4'hb == lineCounter ? frameBuffer_11_39 : _GEN_2811; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2813 = 4'hc == lineCounter ? frameBuffer_12_39 : _GEN_2812; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2814 = 4'hd == lineCounter ? frameBuffer_13_39 : _GEN_2813; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2815 = 4'he == lineCounter ? frameBuffer_14_39 : _GEN_2814; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2818 = 4'h1 == lineCounter ? frameBuffer_1_40 : frameBuffer_0_40; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2819 = 4'h2 == lineCounter ? frameBuffer_2_40 : _GEN_2818; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2820 = 4'h3 == lineCounter ? frameBuffer_3_40 : _GEN_2819; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2821 = 4'h4 == lineCounter ? frameBuffer_4_40 : _GEN_2820; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2822 = 4'h5 == lineCounter ? frameBuffer_5_40 : _GEN_2821; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2823 = 4'h6 == lineCounter ? frameBuffer_6_40 : _GEN_2822; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2824 = 4'h7 == lineCounter ? frameBuffer_7_40 : _GEN_2823; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2825 = 4'h8 == lineCounter ? frameBuffer_8_40 : _GEN_2824; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2826 = 4'h9 == lineCounter ? frameBuffer_9_40 : _GEN_2825; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2827 = 4'ha == lineCounter ? frameBuffer_10_40 : _GEN_2826; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2828 = 4'hb == lineCounter ? frameBuffer_11_40 : _GEN_2827; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2829 = 4'hc == lineCounter ? frameBuffer_12_40 : _GEN_2828; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2830 = 4'hd == lineCounter ? frameBuffer_13_40 : _GEN_2829; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2831 = 4'he == lineCounter ? frameBuffer_14_40 : _GEN_2830; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2834 = 4'h1 == lineCounter ? frameBuffer_1_41 : frameBuffer_0_41; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2835 = 4'h2 == lineCounter ? frameBuffer_2_41 : _GEN_2834; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2836 = 4'h3 == lineCounter ? frameBuffer_3_41 : _GEN_2835; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2837 = 4'h4 == lineCounter ? frameBuffer_4_41 : _GEN_2836; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2838 = 4'h5 == lineCounter ? frameBuffer_5_41 : _GEN_2837; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2839 = 4'h6 == lineCounter ? frameBuffer_6_41 : _GEN_2838; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2840 = 4'h7 == lineCounter ? frameBuffer_7_41 : _GEN_2839; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2841 = 4'h8 == lineCounter ? frameBuffer_8_41 : _GEN_2840; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2842 = 4'h9 == lineCounter ? frameBuffer_9_41 : _GEN_2841; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2843 = 4'ha == lineCounter ? frameBuffer_10_41 : _GEN_2842; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2844 = 4'hb == lineCounter ? frameBuffer_11_41 : _GEN_2843; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2845 = 4'hc == lineCounter ? frameBuffer_12_41 : _GEN_2844; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2846 = 4'hd == lineCounter ? frameBuffer_13_41 : _GEN_2845; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2847 = 4'he == lineCounter ? frameBuffer_14_41 : _GEN_2846; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2850 = 4'h1 == lineCounter ? frameBuffer_1_42 : frameBuffer_0_42; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2851 = 4'h2 == lineCounter ? frameBuffer_2_42 : _GEN_2850; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2852 = 4'h3 == lineCounter ? frameBuffer_3_42 : _GEN_2851; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2853 = 4'h4 == lineCounter ? frameBuffer_4_42 : _GEN_2852; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2854 = 4'h5 == lineCounter ? frameBuffer_5_42 : _GEN_2853; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2855 = 4'h6 == lineCounter ? frameBuffer_6_42 : _GEN_2854; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2856 = 4'h7 == lineCounter ? frameBuffer_7_42 : _GEN_2855; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2857 = 4'h8 == lineCounter ? frameBuffer_8_42 : _GEN_2856; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2858 = 4'h9 == lineCounter ? frameBuffer_9_42 : _GEN_2857; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2859 = 4'ha == lineCounter ? frameBuffer_10_42 : _GEN_2858; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2860 = 4'hb == lineCounter ? frameBuffer_11_42 : _GEN_2859; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2861 = 4'hc == lineCounter ? frameBuffer_12_42 : _GEN_2860; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2862 = 4'hd == lineCounter ? frameBuffer_13_42 : _GEN_2861; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2863 = 4'he == lineCounter ? frameBuffer_14_42 : _GEN_2862; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2866 = 4'h1 == lineCounter ? frameBuffer_1_43 : frameBuffer_0_43; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2867 = 4'h2 == lineCounter ? frameBuffer_2_43 : _GEN_2866; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2868 = 4'h3 == lineCounter ? frameBuffer_3_43 : _GEN_2867; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2869 = 4'h4 == lineCounter ? frameBuffer_4_43 : _GEN_2868; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2870 = 4'h5 == lineCounter ? frameBuffer_5_43 : _GEN_2869; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2871 = 4'h6 == lineCounter ? frameBuffer_6_43 : _GEN_2870; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2872 = 4'h7 == lineCounter ? frameBuffer_7_43 : _GEN_2871; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2873 = 4'h8 == lineCounter ? frameBuffer_8_43 : _GEN_2872; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2874 = 4'h9 == lineCounter ? frameBuffer_9_43 : _GEN_2873; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2875 = 4'ha == lineCounter ? frameBuffer_10_43 : _GEN_2874; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2876 = 4'hb == lineCounter ? frameBuffer_11_43 : _GEN_2875; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2877 = 4'hc == lineCounter ? frameBuffer_12_43 : _GEN_2876; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2878 = 4'hd == lineCounter ? frameBuffer_13_43 : _GEN_2877; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2879 = 4'he == lineCounter ? frameBuffer_14_43 : _GEN_2878; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2882 = 4'h1 == lineCounter ? frameBuffer_1_44 : frameBuffer_0_44; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2883 = 4'h2 == lineCounter ? frameBuffer_2_44 : _GEN_2882; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2884 = 4'h3 == lineCounter ? frameBuffer_3_44 : _GEN_2883; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2885 = 4'h4 == lineCounter ? frameBuffer_4_44 : _GEN_2884; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2886 = 4'h5 == lineCounter ? frameBuffer_5_44 : _GEN_2885; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2887 = 4'h6 == lineCounter ? frameBuffer_6_44 : _GEN_2886; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2888 = 4'h7 == lineCounter ? frameBuffer_7_44 : _GEN_2887; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2889 = 4'h8 == lineCounter ? frameBuffer_8_44 : _GEN_2888; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2890 = 4'h9 == lineCounter ? frameBuffer_9_44 : _GEN_2889; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2891 = 4'ha == lineCounter ? frameBuffer_10_44 : _GEN_2890; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2892 = 4'hb == lineCounter ? frameBuffer_11_44 : _GEN_2891; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2893 = 4'hc == lineCounter ? frameBuffer_12_44 : _GEN_2892; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2894 = 4'hd == lineCounter ? frameBuffer_13_44 : _GEN_2893; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2895 = 4'he == lineCounter ? frameBuffer_14_44 : _GEN_2894; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2898 = 4'h1 == lineCounter ? frameBuffer_1_45 : frameBuffer_0_45; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2899 = 4'h2 == lineCounter ? frameBuffer_2_45 : _GEN_2898; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2900 = 4'h3 == lineCounter ? frameBuffer_3_45 : _GEN_2899; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2901 = 4'h4 == lineCounter ? frameBuffer_4_45 : _GEN_2900; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2902 = 4'h5 == lineCounter ? frameBuffer_5_45 : _GEN_2901; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2903 = 4'h6 == lineCounter ? frameBuffer_6_45 : _GEN_2902; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2904 = 4'h7 == lineCounter ? frameBuffer_7_45 : _GEN_2903; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2905 = 4'h8 == lineCounter ? frameBuffer_8_45 : _GEN_2904; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2906 = 4'h9 == lineCounter ? frameBuffer_9_45 : _GEN_2905; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2907 = 4'ha == lineCounter ? frameBuffer_10_45 : _GEN_2906; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2908 = 4'hb == lineCounter ? frameBuffer_11_45 : _GEN_2907; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2909 = 4'hc == lineCounter ? frameBuffer_12_45 : _GEN_2908; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2910 = 4'hd == lineCounter ? frameBuffer_13_45 : _GEN_2909; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2911 = 4'he == lineCounter ? frameBuffer_14_45 : _GEN_2910; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2914 = 4'h1 == lineCounter ? frameBuffer_1_46 : frameBuffer_0_46; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2915 = 4'h2 == lineCounter ? frameBuffer_2_46 : _GEN_2914; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2916 = 4'h3 == lineCounter ? frameBuffer_3_46 : _GEN_2915; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2917 = 4'h4 == lineCounter ? frameBuffer_4_46 : _GEN_2916; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2918 = 4'h5 == lineCounter ? frameBuffer_5_46 : _GEN_2917; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2919 = 4'h6 == lineCounter ? frameBuffer_6_46 : _GEN_2918; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2920 = 4'h7 == lineCounter ? frameBuffer_7_46 : _GEN_2919; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2921 = 4'h8 == lineCounter ? frameBuffer_8_46 : _GEN_2920; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2922 = 4'h9 == lineCounter ? frameBuffer_9_46 : _GEN_2921; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2923 = 4'ha == lineCounter ? frameBuffer_10_46 : _GEN_2922; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2924 = 4'hb == lineCounter ? frameBuffer_11_46 : _GEN_2923; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2925 = 4'hc == lineCounter ? frameBuffer_12_46 : _GEN_2924; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2926 = 4'hd == lineCounter ? frameBuffer_13_46 : _GEN_2925; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2927 = 4'he == lineCounter ? frameBuffer_14_46 : _GEN_2926; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2930 = 4'h1 == lineCounter ? frameBuffer_1_47 : frameBuffer_0_47; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2931 = 4'h2 == lineCounter ? frameBuffer_2_47 : _GEN_2930; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2932 = 4'h3 == lineCounter ? frameBuffer_3_47 : _GEN_2931; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2933 = 4'h4 == lineCounter ? frameBuffer_4_47 : _GEN_2932; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2934 = 4'h5 == lineCounter ? frameBuffer_5_47 : _GEN_2933; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2935 = 4'h6 == lineCounter ? frameBuffer_6_47 : _GEN_2934; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2936 = 4'h7 == lineCounter ? frameBuffer_7_47 : _GEN_2935; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2937 = 4'h8 == lineCounter ? frameBuffer_8_47 : _GEN_2936; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2938 = 4'h9 == lineCounter ? frameBuffer_9_47 : _GEN_2937; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2939 = 4'ha == lineCounter ? frameBuffer_10_47 : _GEN_2938; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2940 = 4'hb == lineCounter ? frameBuffer_11_47 : _GEN_2939; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2941 = 4'hc == lineCounter ? frameBuffer_12_47 : _GEN_2940; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2942 = 4'hd == lineCounter ? frameBuffer_13_47 : _GEN_2941; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2943 = 4'he == lineCounter ? frameBuffer_14_47 : _GEN_2942; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2946 = 4'h1 == lineCounter ? frameBuffer_1_48 : frameBuffer_0_48; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2947 = 4'h2 == lineCounter ? frameBuffer_2_48 : _GEN_2946; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2948 = 4'h3 == lineCounter ? frameBuffer_3_48 : _GEN_2947; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2949 = 4'h4 == lineCounter ? frameBuffer_4_48 : _GEN_2948; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2950 = 4'h5 == lineCounter ? frameBuffer_5_48 : _GEN_2949; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2951 = 4'h6 == lineCounter ? frameBuffer_6_48 : _GEN_2950; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2952 = 4'h7 == lineCounter ? frameBuffer_7_48 : _GEN_2951; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2953 = 4'h8 == lineCounter ? frameBuffer_8_48 : _GEN_2952; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2954 = 4'h9 == lineCounter ? frameBuffer_9_48 : _GEN_2953; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2955 = 4'ha == lineCounter ? frameBuffer_10_48 : _GEN_2954; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2956 = 4'hb == lineCounter ? frameBuffer_11_48 : _GEN_2955; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2957 = 4'hc == lineCounter ? frameBuffer_12_48 : _GEN_2956; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2958 = 4'hd == lineCounter ? frameBuffer_13_48 : _GEN_2957; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2959 = 4'he == lineCounter ? frameBuffer_14_48 : _GEN_2958; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2962 = 4'h1 == lineCounter ? frameBuffer_1_49 : frameBuffer_0_49; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2963 = 4'h2 == lineCounter ? frameBuffer_2_49 : _GEN_2962; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2964 = 4'h3 == lineCounter ? frameBuffer_3_49 : _GEN_2963; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2965 = 4'h4 == lineCounter ? frameBuffer_4_49 : _GEN_2964; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2966 = 4'h5 == lineCounter ? frameBuffer_5_49 : _GEN_2965; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2967 = 4'h6 == lineCounter ? frameBuffer_6_49 : _GEN_2966; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2968 = 4'h7 == lineCounter ? frameBuffer_7_49 : _GEN_2967; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2969 = 4'h8 == lineCounter ? frameBuffer_8_49 : _GEN_2968; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2970 = 4'h9 == lineCounter ? frameBuffer_9_49 : _GEN_2969; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2971 = 4'ha == lineCounter ? frameBuffer_10_49 : _GEN_2970; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2972 = 4'hb == lineCounter ? frameBuffer_11_49 : _GEN_2971; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2973 = 4'hc == lineCounter ? frameBuffer_12_49 : _GEN_2972; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2974 = 4'hd == lineCounter ? frameBuffer_13_49 : _GEN_2973; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2975 = 4'he == lineCounter ? frameBuffer_14_49 : _GEN_2974; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2978 = 4'h1 == lineCounter ? frameBuffer_1_50 : frameBuffer_0_50; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2979 = 4'h2 == lineCounter ? frameBuffer_2_50 : _GEN_2978; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2980 = 4'h3 == lineCounter ? frameBuffer_3_50 : _GEN_2979; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2981 = 4'h4 == lineCounter ? frameBuffer_4_50 : _GEN_2980; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2982 = 4'h5 == lineCounter ? frameBuffer_5_50 : _GEN_2981; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2983 = 4'h6 == lineCounter ? frameBuffer_6_50 : _GEN_2982; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2984 = 4'h7 == lineCounter ? frameBuffer_7_50 : _GEN_2983; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2985 = 4'h8 == lineCounter ? frameBuffer_8_50 : _GEN_2984; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2986 = 4'h9 == lineCounter ? frameBuffer_9_50 : _GEN_2985; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2987 = 4'ha == lineCounter ? frameBuffer_10_50 : _GEN_2986; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2988 = 4'hb == lineCounter ? frameBuffer_11_50 : _GEN_2987; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2989 = 4'hc == lineCounter ? frameBuffer_12_50 : _GEN_2988; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2990 = 4'hd == lineCounter ? frameBuffer_13_50 : _GEN_2989; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2991 = 4'he == lineCounter ? frameBuffer_14_50 : _GEN_2990; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2994 = 4'h1 == lineCounter ? frameBuffer_1_51 : frameBuffer_0_51; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2995 = 4'h2 == lineCounter ? frameBuffer_2_51 : _GEN_2994; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2996 = 4'h3 == lineCounter ? frameBuffer_3_51 : _GEN_2995; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2997 = 4'h4 == lineCounter ? frameBuffer_4_51 : _GEN_2996; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2998 = 4'h5 == lineCounter ? frameBuffer_5_51 : _GEN_2997; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_2999 = 4'h6 == lineCounter ? frameBuffer_6_51 : _GEN_2998; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3000 = 4'h7 == lineCounter ? frameBuffer_7_51 : _GEN_2999; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3001 = 4'h8 == lineCounter ? frameBuffer_8_51 : _GEN_3000; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3002 = 4'h9 == lineCounter ? frameBuffer_9_51 : _GEN_3001; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3003 = 4'ha == lineCounter ? frameBuffer_10_51 : _GEN_3002; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3004 = 4'hb == lineCounter ? frameBuffer_11_51 : _GEN_3003; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3005 = 4'hc == lineCounter ? frameBuffer_12_51 : _GEN_3004; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3006 = 4'hd == lineCounter ? frameBuffer_13_51 : _GEN_3005; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3007 = 4'he == lineCounter ? frameBuffer_14_51 : _GEN_3006; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3010 = 4'h1 == lineCounter ? frameBuffer_1_52 : frameBuffer_0_52; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3011 = 4'h2 == lineCounter ? frameBuffer_2_52 : _GEN_3010; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3012 = 4'h3 == lineCounter ? frameBuffer_3_52 : _GEN_3011; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3013 = 4'h4 == lineCounter ? frameBuffer_4_52 : _GEN_3012; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3014 = 4'h5 == lineCounter ? frameBuffer_5_52 : _GEN_3013; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3015 = 4'h6 == lineCounter ? frameBuffer_6_52 : _GEN_3014; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3016 = 4'h7 == lineCounter ? frameBuffer_7_52 : _GEN_3015; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3017 = 4'h8 == lineCounter ? frameBuffer_8_52 : _GEN_3016; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3018 = 4'h9 == lineCounter ? frameBuffer_9_52 : _GEN_3017; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3019 = 4'ha == lineCounter ? frameBuffer_10_52 : _GEN_3018; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3020 = 4'hb == lineCounter ? frameBuffer_11_52 : _GEN_3019; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3021 = 4'hc == lineCounter ? frameBuffer_12_52 : _GEN_3020; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3022 = 4'hd == lineCounter ? frameBuffer_13_52 : _GEN_3021; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3023 = 4'he == lineCounter ? frameBuffer_14_52 : _GEN_3022; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3026 = 4'h1 == lineCounter ? frameBuffer_1_53 : frameBuffer_0_53; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3027 = 4'h2 == lineCounter ? frameBuffer_2_53 : _GEN_3026; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3028 = 4'h3 == lineCounter ? frameBuffer_3_53 : _GEN_3027; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3029 = 4'h4 == lineCounter ? frameBuffer_4_53 : _GEN_3028; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3030 = 4'h5 == lineCounter ? frameBuffer_5_53 : _GEN_3029; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3031 = 4'h6 == lineCounter ? frameBuffer_6_53 : _GEN_3030; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3032 = 4'h7 == lineCounter ? frameBuffer_7_53 : _GEN_3031; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3033 = 4'h8 == lineCounter ? frameBuffer_8_53 : _GEN_3032; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3034 = 4'h9 == lineCounter ? frameBuffer_9_53 : _GEN_3033; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3035 = 4'ha == lineCounter ? frameBuffer_10_53 : _GEN_3034; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3036 = 4'hb == lineCounter ? frameBuffer_11_53 : _GEN_3035; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3037 = 4'hc == lineCounter ? frameBuffer_12_53 : _GEN_3036; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3038 = 4'hd == lineCounter ? frameBuffer_13_53 : _GEN_3037; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3039 = 4'he == lineCounter ? frameBuffer_14_53 : _GEN_3038; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3042 = 4'h1 == lineCounter ? frameBuffer_1_54 : frameBuffer_0_54; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3043 = 4'h2 == lineCounter ? frameBuffer_2_54 : _GEN_3042; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3044 = 4'h3 == lineCounter ? frameBuffer_3_54 : _GEN_3043; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3045 = 4'h4 == lineCounter ? frameBuffer_4_54 : _GEN_3044; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3046 = 4'h5 == lineCounter ? frameBuffer_5_54 : _GEN_3045; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3047 = 4'h6 == lineCounter ? frameBuffer_6_54 : _GEN_3046; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3048 = 4'h7 == lineCounter ? frameBuffer_7_54 : _GEN_3047; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3049 = 4'h8 == lineCounter ? frameBuffer_8_54 : _GEN_3048; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3050 = 4'h9 == lineCounter ? frameBuffer_9_54 : _GEN_3049; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3051 = 4'ha == lineCounter ? frameBuffer_10_54 : _GEN_3050; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3052 = 4'hb == lineCounter ? frameBuffer_11_54 : _GEN_3051; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3053 = 4'hc == lineCounter ? frameBuffer_12_54 : _GEN_3052; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3054 = 4'hd == lineCounter ? frameBuffer_13_54 : _GEN_3053; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3055 = 4'he == lineCounter ? frameBuffer_14_54 : _GEN_3054; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3058 = 4'h1 == lineCounter ? frameBuffer_1_55 : frameBuffer_0_55; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3059 = 4'h2 == lineCounter ? frameBuffer_2_55 : _GEN_3058; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3060 = 4'h3 == lineCounter ? frameBuffer_3_55 : _GEN_3059; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3061 = 4'h4 == lineCounter ? frameBuffer_4_55 : _GEN_3060; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3062 = 4'h5 == lineCounter ? frameBuffer_5_55 : _GEN_3061; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3063 = 4'h6 == lineCounter ? frameBuffer_6_55 : _GEN_3062; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3064 = 4'h7 == lineCounter ? frameBuffer_7_55 : _GEN_3063; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3065 = 4'h8 == lineCounter ? frameBuffer_8_55 : _GEN_3064; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3066 = 4'h9 == lineCounter ? frameBuffer_9_55 : _GEN_3065; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3067 = 4'ha == lineCounter ? frameBuffer_10_55 : _GEN_3066; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3068 = 4'hb == lineCounter ? frameBuffer_11_55 : _GEN_3067; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3069 = 4'hc == lineCounter ? frameBuffer_12_55 : _GEN_3068; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3070 = 4'hd == lineCounter ? frameBuffer_13_55 : _GEN_3069; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3071 = 4'he == lineCounter ? frameBuffer_14_55 : _GEN_3070; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3074 = 4'h1 == lineCounter ? frameBuffer_1_56 : frameBuffer_0_56; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3075 = 4'h2 == lineCounter ? frameBuffer_2_56 : _GEN_3074; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3076 = 4'h3 == lineCounter ? frameBuffer_3_56 : _GEN_3075; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3077 = 4'h4 == lineCounter ? frameBuffer_4_56 : _GEN_3076; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3078 = 4'h5 == lineCounter ? frameBuffer_5_56 : _GEN_3077; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3079 = 4'h6 == lineCounter ? frameBuffer_6_56 : _GEN_3078; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3080 = 4'h7 == lineCounter ? frameBuffer_7_56 : _GEN_3079; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3081 = 4'h8 == lineCounter ? frameBuffer_8_56 : _GEN_3080; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3082 = 4'h9 == lineCounter ? frameBuffer_9_56 : _GEN_3081; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3083 = 4'ha == lineCounter ? frameBuffer_10_56 : _GEN_3082; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3084 = 4'hb == lineCounter ? frameBuffer_11_56 : _GEN_3083; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3085 = 4'hc == lineCounter ? frameBuffer_12_56 : _GEN_3084; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3086 = 4'hd == lineCounter ? frameBuffer_13_56 : _GEN_3085; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3087 = 4'he == lineCounter ? frameBuffer_14_56 : _GEN_3086; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3090 = 4'h1 == lineCounter ? frameBuffer_1_57 : frameBuffer_0_57; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3091 = 4'h2 == lineCounter ? frameBuffer_2_57 : _GEN_3090; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3092 = 4'h3 == lineCounter ? frameBuffer_3_57 : _GEN_3091; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3093 = 4'h4 == lineCounter ? frameBuffer_4_57 : _GEN_3092; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3094 = 4'h5 == lineCounter ? frameBuffer_5_57 : _GEN_3093; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3095 = 4'h6 == lineCounter ? frameBuffer_6_57 : _GEN_3094; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3096 = 4'h7 == lineCounter ? frameBuffer_7_57 : _GEN_3095; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3097 = 4'h8 == lineCounter ? frameBuffer_8_57 : _GEN_3096; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3098 = 4'h9 == lineCounter ? frameBuffer_9_57 : _GEN_3097; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3099 = 4'ha == lineCounter ? frameBuffer_10_57 : _GEN_3098; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3100 = 4'hb == lineCounter ? frameBuffer_11_57 : _GEN_3099; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3101 = 4'hc == lineCounter ? frameBuffer_12_57 : _GEN_3100; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3102 = 4'hd == lineCounter ? frameBuffer_13_57 : _GEN_3101; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3103 = 4'he == lineCounter ? frameBuffer_14_57 : _GEN_3102; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3106 = 4'h1 == lineCounter ? frameBuffer_1_58 : frameBuffer_0_58; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3107 = 4'h2 == lineCounter ? frameBuffer_2_58 : _GEN_3106; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3108 = 4'h3 == lineCounter ? frameBuffer_3_58 : _GEN_3107; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3109 = 4'h4 == lineCounter ? frameBuffer_4_58 : _GEN_3108; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3110 = 4'h5 == lineCounter ? frameBuffer_5_58 : _GEN_3109; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3111 = 4'h6 == lineCounter ? frameBuffer_6_58 : _GEN_3110; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3112 = 4'h7 == lineCounter ? frameBuffer_7_58 : _GEN_3111; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3113 = 4'h8 == lineCounter ? frameBuffer_8_58 : _GEN_3112; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3114 = 4'h9 == lineCounter ? frameBuffer_9_58 : _GEN_3113; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3115 = 4'ha == lineCounter ? frameBuffer_10_58 : _GEN_3114; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3116 = 4'hb == lineCounter ? frameBuffer_11_58 : _GEN_3115; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3117 = 4'hc == lineCounter ? frameBuffer_12_58 : _GEN_3116; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3118 = 4'hd == lineCounter ? frameBuffer_13_58 : _GEN_3117; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3119 = 4'he == lineCounter ? frameBuffer_14_58 : _GEN_3118; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3122 = 4'h1 == lineCounter ? frameBuffer_1_59 : frameBuffer_0_59; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3123 = 4'h2 == lineCounter ? frameBuffer_2_59 : _GEN_3122; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3124 = 4'h3 == lineCounter ? frameBuffer_3_59 : _GEN_3123; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3125 = 4'h4 == lineCounter ? frameBuffer_4_59 : _GEN_3124; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3126 = 4'h5 == lineCounter ? frameBuffer_5_59 : _GEN_3125; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3127 = 4'h6 == lineCounter ? frameBuffer_6_59 : _GEN_3126; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3128 = 4'h7 == lineCounter ? frameBuffer_7_59 : _GEN_3127; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3129 = 4'h8 == lineCounter ? frameBuffer_8_59 : _GEN_3128; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3130 = 4'h9 == lineCounter ? frameBuffer_9_59 : _GEN_3129; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3131 = 4'ha == lineCounter ? frameBuffer_10_59 : _GEN_3130; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3132 = 4'hb == lineCounter ? frameBuffer_11_59 : _GEN_3131; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3133 = 4'hc == lineCounter ? frameBuffer_12_59 : _GEN_3132; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3134 = 4'hd == lineCounter ? frameBuffer_13_59 : _GEN_3133; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3135 = 4'he == lineCounter ? frameBuffer_14_59 : _GEN_3134; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3138 = 4'h1 == lineCounter ? frameBuffer_1_60 : frameBuffer_0_60; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3139 = 4'h2 == lineCounter ? frameBuffer_2_60 : _GEN_3138; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3140 = 4'h3 == lineCounter ? frameBuffer_3_60 : _GEN_3139; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3141 = 4'h4 == lineCounter ? frameBuffer_4_60 : _GEN_3140; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3142 = 4'h5 == lineCounter ? frameBuffer_5_60 : _GEN_3141; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3143 = 4'h6 == lineCounter ? frameBuffer_6_60 : _GEN_3142; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3144 = 4'h7 == lineCounter ? frameBuffer_7_60 : _GEN_3143; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3145 = 4'h8 == lineCounter ? frameBuffer_8_60 : _GEN_3144; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3146 = 4'h9 == lineCounter ? frameBuffer_9_60 : _GEN_3145; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3147 = 4'ha == lineCounter ? frameBuffer_10_60 : _GEN_3146; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3148 = 4'hb == lineCounter ? frameBuffer_11_60 : _GEN_3147; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3149 = 4'hc == lineCounter ? frameBuffer_12_60 : _GEN_3148; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3150 = 4'hd == lineCounter ? frameBuffer_13_60 : _GEN_3149; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3151 = 4'he == lineCounter ? frameBuffer_14_60 : _GEN_3150; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3154 = 4'h1 == lineCounter ? frameBuffer_1_61 : frameBuffer_0_61; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3155 = 4'h2 == lineCounter ? frameBuffer_2_61 : _GEN_3154; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3156 = 4'h3 == lineCounter ? frameBuffer_3_61 : _GEN_3155; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3157 = 4'h4 == lineCounter ? frameBuffer_4_61 : _GEN_3156; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3158 = 4'h5 == lineCounter ? frameBuffer_5_61 : _GEN_3157; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3159 = 4'h6 == lineCounter ? frameBuffer_6_61 : _GEN_3158; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3160 = 4'h7 == lineCounter ? frameBuffer_7_61 : _GEN_3159; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3161 = 4'h8 == lineCounter ? frameBuffer_8_61 : _GEN_3160; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3162 = 4'h9 == lineCounter ? frameBuffer_9_61 : _GEN_3161; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3163 = 4'ha == lineCounter ? frameBuffer_10_61 : _GEN_3162; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3164 = 4'hb == lineCounter ? frameBuffer_11_61 : _GEN_3163; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3165 = 4'hc == lineCounter ? frameBuffer_12_61 : _GEN_3164; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3166 = 4'hd == lineCounter ? frameBuffer_13_61 : _GEN_3165; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3167 = 4'he == lineCounter ? frameBuffer_14_61 : _GEN_3166; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3170 = 4'h1 == lineCounter ? frameBuffer_1_62 : frameBuffer_0_62; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3171 = 4'h2 == lineCounter ? frameBuffer_2_62 : _GEN_3170; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3172 = 4'h3 == lineCounter ? frameBuffer_3_62 : _GEN_3171; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3173 = 4'h4 == lineCounter ? frameBuffer_4_62 : _GEN_3172; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3174 = 4'h5 == lineCounter ? frameBuffer_5_62 : _GEN_3173; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3175 = 4'h6 == lineCounter ? frameBuffer_6_62 : _GEN_3174; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3176 = 4'h7 == lineCounter ? frameBuffer_7_62 : _GEN_3175; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3177 = 4'h8 == lineCounter ? frameBuffer_8_62 : _GEN_3176; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3178 = 4'h9 == lineCounter ? frameBuffer_9_62 : _GEN_3177; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3179 = 4'ha == lineCounter ? frameBuffer_10_62 : _GEN_3178; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3180 = 4'hb == lineCounter ? frameBuffer_11_62 : _GEN_3179; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3181 = 4'hc == lineCounter ? frameBuffer_12_62 : _GEN_3180; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3182 = 4'hd == lineCounter ? frameBuffer_13_62 : _GEN_3181; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3183 = 4'he == lineCounter ? frameBuffer_14_62 : _GEN_3182; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3186 = 4'h1 == lineCounter ? frameBuffer_1_63 : frameBuffer_0_63; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3187 = 4'h2 == lineCounter ? frameBuffer_2_63 : _GEN_3186; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3188 = 4'h3 == lineCounter ? frameBuffer_3_63 : _GEN_3187; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3189 = 4'h4 == lineCounter ? frameBuffer_4_63 : _GEN_3188; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3190 = 4'h5 == lineCounter ? frameBuffer_5_63 : _GEN_3189; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3191 = 4'h6 == lineCounter ? frameBuffer_6_63 : _GEN_3190; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3192 = 4'h7 == lineCounter ? frameBuffer_7_63 : _GEN_3191; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3193 = 4'h8 == lineCounter ? frameBuffer_8_63 : _GEN_3192; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3194 = 4'h9 == lineCounter ? frameBuffer_9_63 : _GEN_3193; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3195 = 4'ha == lineCounter ? frameBuffer_10_63 : _GEN_3194; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3196 = 4'hb == lineCounter ? frameBuffer_11_63 : _GEN_3195; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3197 = 4'hc == lineCounter ? frameBuffer_12_63 : _GEN_3196; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3198 = 4'hd == lineCounter ? frameBuffer_13_63 : _GEN_3197; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3199 = 4'he == lineCounter ? frameBuffer_14_63 : _GEN_3198; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3202 = 4'h1 == lineCounter ? frameBuffer_1_64 : frameBuffer_0_64; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3203 = 4'h2 == lineCounter ? frameBuffer_2_64 : _GEN_3202; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3204 = 4'h3 == lineCounter ? frameBuffer_3_64 : _GEN_3203; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3205 = 4'h4 == lineCounter ? frameBuffer_4_64 : _GEN_3204; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3206 = 4'h5 == lineCounter ? frameBuffer_5_64 : _GEN_3205; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3207 = 4'h6 == lineCounter ? frameBuffer_6_64 : _GEN_3206; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3208 = 4'h7 == lineCounter ? frameBuffer_7_64 : _GEN_3207; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3209 = 4'h8 == lineCounter ? frameBuffer_8_64 : _GEN_3208; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3210 = 4'h9 == lineCounter ? frameBuffer_9_64 : _GEN_3209; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3211 = 4'ha == lineCounter ? frameBuffer_10_64 : _GEN_3210; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3212 = 4'hb == lineCounter ? frameBuffer_11_64 : _GEN_3211; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3213 = 4'hc == lineCounter ? frameBuffer_12_64 : _GEN_3212; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3214 = 4'hd == lineCounter ? frameBuffer_13_64 : _GEN_3213; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3215 = 4'he == lineCounter ? frameBuffer_14_64 : _GEN_3214; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3218 = 4'h1 == lineCounter ? frameBuffer_1_65 : frameBuffer_0_65; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3219 = 4'h2 == lineCounter ? frameBuffer_2_65 : _GEN_3218; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3220 = 4'h3 == lineCounter ? frameBuffer_3_65 : _GEN_3219; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3221 = 4'h4 == lineCounter ? frameBuffer_4_65 : _GEN_3220; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3222 = 4'h5 == lineCounter ? frameBuffer_5_65 : _GEN_3221; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3223 = 4'h6 == lineCounter ? frameBuffer_6_65 : _GEN_3222; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3224 = 4'h7 == lineCounter ? frameBuffer_7_65 : _GEN_3223; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3225 = 4'h8 == lineCounter ? frameBuffer_8_65 : _GEN_3224; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3226 = 4'h9 == lineCounter ? frameBuffer_9_65 : _GEN_3225; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3227 = 4'ha == lineCounter ? frameBuffer_10_65 : _GEN_3226; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3228 = 4'hb == lineCounter ? frameBuffer_11_65 : _GEN_3227; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3229 = 4'hc == lineCounter ? frameBuffer_12_65 : _GEN_3228; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3230 = 4'hd == lineCounter ? frameBuffer_13_65 : _GEN_3229; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3231 = 4'he == lineCounter ? frameBuffer_14_65 : _GEN_3230; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3234 = 4'h1 == lineCounter ? frameBuffer_1_66 : frameBuffer_0_66; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3235 = 4'h2 == lineCounter ? frameBuffer_2_66 : _GEN_3234; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3236 = 4'h3 == lineCounter ? frameBuffer_3_66 : _GEN_3235; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3237 = 4'h4 == lineCounter ? frameBuffer_4_66 : _GEN_3236; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3238 = 4'h5 == lineCounter ? frameBuffer_5_66 : _GEN_3237; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3239 = 4'h6 == lineCounter ? frameBuffer_6_66 : _GEN_3238; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3240 = 4'h7 == lineCounter ? frameBuffer_7_66 : _GEN_3239; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3241 = 4'h8 == lineCounter ? frameBuffer_8_66 : _GEN_3240; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3242 = 4'h9 == lineCounter ? frameBuffer_9_66 : _GEN_3241; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3243 = 4'ha == lineCounter ? frameBuffer_10_66 : _GEN_3242; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3244 = 4'hb == lineCounter ? frameBuffer_11_66 : _GEN_3243; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3245 = 4'hc == lineCounter ? frameBuffer_12_66 : _GEN_3244; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3246 = 4'hd == lineCounter ? frameBuffer_13_66 : _GEN_3245; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3247 = 4'he == lineCounter ? frameBuffer_14_66 : _GEN_3246; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3250 = 4'h1 == lineCounter ? frameBuffer_1_67 : frameBuffer_0_67; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3251 = 4'h2 == lineCounter ? frameBuffer_2_67 : _GEN_3250; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3252 = 4'h3 == lineCounter ? frameBuffer_3_67 : _GEN_3251; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3253 = 4'h4 == lineCounter ? frameBuffer_4_67 : _GEN_3252; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3254 = 4'h5 == lineCounter ? frameBuffer_5_67 : _GEN_3253; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3255 = 4'h6 == lineCounter ? frameBuffer_6_67 : _GEN_3254; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3256 = 4'h7 == lineCounter ? frameBuffer_7_67 : _GEN_3255; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3257 = 4'h8 == lineCounter ? frameBuffer_8_67 : _GEN_3256; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3258 = 4'h9 == lineCounter ? frameBuffer_9_67 : _GEN_3257; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3259 = 4'ha == lineCounter ? frameBuffer_10_67 : _GEN_3258; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3260 = 4'hb == lineCounter ? frameBuffer_11_67 : _GEN_3259; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3261 = 4'hc == lineCounter ? frameBuffer_12_67 : _GEN_3260; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3262 = 4'hd == lineCounter ? frameBuffer_13_67 : _GEN_3261; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3263 = 4'he == lineCounter ? frameBuffer_14_67 : _GEN_3262; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3266 = 4'h1 == lineCounter ? frameBuffer_1_68 : frameBuffer_0_68; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3267 = 4'h2 == lineCounter ? frameBuffer_2_68 : _GEN_3266; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3268 = 4'h3 == lineCounter ? frameBuffer_3_68 : _GEN_3267; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3269 = 4'h4 == lineCounter ? frameBuffer_4_68 : _GEN_3268; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3270 = 4'h5 == lineCounter ? frameBuffer_5_68 : _GEN_3269; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3271 = 4'h6 == lineCounter ? frameBuffer_6_68 : _GEN_3270; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3272 = 4'h7 == lineCounter ? frameBuffer_7_68 : _GEN_3271; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3273 = 4'h8 == lineCounter ? frameBuffer_8_68 : _GEN_3272; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3274 = 4'h9 == lineCounter ? frameBuffer_9_68 : _GEN_3273; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3275 = 4'ha == lineCounter ? frameBuffer_10_68 : _GEN_3274; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3276 = 4'hb == lineCounter ? frameBuffer_11_68 : _GEN_3275; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3277 = 4'hc == lineCounter ? frameBuffer_12_68 : _GEN_3276; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3278 = 4'hd == lineCounter ? frameBuffer_13_68 : _GEN_3277; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3279 = 4'he == lineCounter ? frameBuffer_14_68 : _GEN_3278; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3282 = 4'h1 == lineCounter ? frameBuffer_1_69 : frameBuffer_0_69; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3283 = 4'h2 == lineCounter ? frameBuffer_2_69 : _GEN_3282; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3284 = 4'h3 == lineCounter ? frameBuffer_3_69 : _GEN_3283; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3285 = 4'h4 == lineCounter ? frameBuffer_4_69 : _GEN_3284; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3286 = 4'h5 == lineCounter ? frameBuffer_5_69 : _GEN_3285; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3287 = 4'h6 == lineCounter ? frameBuffer_6_69 : _GEN_3286; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3288 = 4'h7 == lineCounter ? frameBuffer_7_69 : _GEN_3287; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3289 = 4'h8 == lineCounter ? frameBuffer_8_69 : _GEN_3288; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3290 = 4'h9 == lineCounter ? frameBuffer_9_69 : _GEN_3289; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3291 = 4'ha == lineCounter ? frameBuffer_10_69 : _GEN_3290; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3292 = 4'hb == lineCounter ? frameBuffer_11_69 : _GEN_3291; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3293 = 4'hc == lineCounter ? frameBuffer_12_69 : _GEN_3292; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3294 = 4'hd == lineCounter ? frameBuffer_13_69 : _GEN_3293; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3295 = 4'he == lineCounter ? frameBuffer_14_69 : _GEN_3294; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3298 = 4'h1 == lineCounter ? frameBuffer_1_70 : frameBuffer_0_70; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3299 = 4'h2 == lineCounter ? frameBuffer_2_70 : _GEN_3298; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3300 = 4'h3 == lineCounter ? frameBuffer_3_70 : _GEN_3299; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3301 = 4'h4 == lineCounter ? frameBuffer_4_70 : _GEN_3300; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3302 = 4'h5 == lineCounter ? frameBuffer_5_70 : _GEN_3301; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3303 = 4'h6 == lineCounter ? frameBuffer_6_70 : _GEN_3302; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3304 = 4'h7 == lineCounter ? frameBuffer_7_70 : _GEN_3303; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3305 = 4'h8 == lineCounter ? frameBuffer_8_70 : _GEN_3304; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3306 = 4'h9 == lineCounter ? frameBuffer_9_70 : _GEN_3305; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3307 = 4'ha == lineCounter ? frameBuffer_10_70 : _GEN_3306; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3308 = 4'hb == lineCounter ? frameBuffer_11_70 : _GEN_3307; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3309 = 4'hc == lineCounter ? frameBuffer_12_70 : _GEN_3308; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3310 = 4'hd == lineCounter ? frameBuffer_13_70 : _GEN_3309; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3311 = 4'he == lineCounter ? frameBuffer_14_70 : _GEN_3310; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3314 = 4'h1 == lineCounter ? frameBuffer_1_71 : frameBuffer_0_71; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3315 = 4'h2 == lineCounter ? frameBuffer_2_71 : _GEN_3314; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3316 = 4'h3 == lineCounter ? frameBuffer_3_71 : _GEN_3315; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3317 = 4'h4 == lineCounter ? frameBuffer_4_71 : _GEN_3316; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3318 = 4'h5 == lineCounter ? frameBuffer_5_71 : _GEN_3317; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3319 = 4'h6 == lineCounter ? frameBuffer_6_71 : _GEN_3318; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3320 = 4'h7 == lineCounter ? frameBuffer_7_71 : _GEN_3319; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3321 = 4'h8 == lineCounter ? frameBuffer_8_71 : _GEN_3320; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3322 = 4'h9 == lineCounter ? frameBuffer_9_71 : _GEN_3321; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3323 = 4'ha == lineCounter ? frameBuffer_10_71 : _GEN_3322; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3324 = 4'hb == lineCounter ? frameBuffer_11_71 : _GEN_3323; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3325 = 4'hc == lineCounter ? frameBuffer_12_71 : _GEN_3324; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3326 = 4'hd == lineCounter ? frameBuffer_13_71 : _GEN_3325; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3327 = 4'he == lineCounter ? frameBuffer_14_71 : _GEN_3326; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3330 = 4'h1 == lineCounter ? frameBuffer_1_72 : frameBuffer_0_72; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3331 = 4'h2 == lineCounter ? frameBuffer_2_72 : _GEN_3330; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3332 = 4'h3 == lineCounter ? frameBuffer_3_72 : _GEN_3331; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3333 = 4'h4 == lineCounter ? frameBuffer_4_72 : _GEN_3332; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3334 = 4'h5 == lineCounter ? frameBuffer_5_72 : _GEN_3333; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3335 = 4'h6 == lineCounter ? frameBuffer_6_72 : _GEN_3334; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3336 = 4'h7 == lineCounter ? frameBuffer_7_72 : _GEN_3335; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3337 = 4'h8 == lineCounter ? frameBuffer_8_72 : _GEN_3336; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3338 = 4'h9 == lineCounter ? frameBuffer_9_72 : _GEN_3337; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3339 = 4'ha == lineCounter ? frameBuffer_10_72 : _GEN_3338; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3340 = 4'hb == lineCounter ? frameBuffer_11_72 : _GEN_3339; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3341 = 4'hc == lineCounter ? frameBuffer_12_72 : _GEN_3340; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3342 = 4'hd == lineCounter ? frameBuffer_13_72 : _GEN_3341; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3343 = 4'he == lineCounter ? frameBuffer_14_72 : _GEN_3342; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3346 = 4'h1 == lineCounter ? frameBuffer_1_73 : frameBuffer_0_73; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3347 = 4'h2 == lineCounter ? frameBuffer_2_73 : _GEN_3346; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3348 = 4'h3 == lineCounter ? frameBuffer_3_73 : _GEN_3347; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3349 = 4'h4 == lineCounter ? frameBuffer_4_73 : _GEN_3348; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3350 = 4'h5 == lineCounter ? frameBuffer_5_73 : _GEN_3349; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3351 = 4'h6 == lineCounter ? frameBuffer_6_73 : _GEN_3350; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3352 = 4'h7 == lineCounter ? frameBuffer_7_73 : _GEN_3351; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3353 = 4'h8 == lineCounter ? frameBuffer_8_73 : _GEN_3352; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3354 = 4'h9 == lineCounter ? frameBuffer_9_73 : _GEN_3353; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3355 = 4'ha == lineCounter ? frameBuffer_10_73 : _GEN_3354; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3356 = 4'hb == lineCounter ? frameBuffer_11_73 : _GEN_3355; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3357 = 4'hc == lineCounter ? frameBuffer_12_73 : _GEN_3356; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3358 = 4'hd == lineCounter ? frameBuffer_13_73 : _GEN_3357; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3359 = 4'he == lineCounter ? frameBuffer_14_73 : _GEN_3358; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3362 = 4'h1 == lineCounter ? frameBuffer_1_74 : frameBuffer_0_74; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3363 = 4'h2 == lineCounter ? frameBuffer_2_74 : _GEN_3362; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3364 = 4'h3 == lineCounter ? frameBuffer_3_74 : _GEN_3363; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3365 = 4'h4 == lineCounter ? frameBuffer_4_74 : _GEN_3364; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3366 = 4'h5 == lineCounter ? frameBuffer_5_74 : _GEN_3365; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3367 = 4'h6 == lineCounter ? frameBuffer_6_74 : _GEN_3366; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3368 = 4'h7 == lineCounter ? frameBuffer_7_74 : _GEN_3367; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3369 = 4'h8 == lineCounter ? frameBuffer_8_74 : _GEN_3368; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3370 = 4'h9 == lineCounter ? frameBuffer_9_74 : _GEN_3369; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3371 = 4'ha == lineCounter ? frameBuffer_10_74 : _GEN_3370; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3372 = 4'hb == lineCounter ? frameBuffer_11_74 : _GEN_3371; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3373 = 4'hc == lineCounter ? frameBuffer_12_74 : _GEN_3372; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3374 = 4'hd == lineCounter ? frameBuffer_13_74 : _GEN_3373; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3375 = 4'he == lineCounter ? frameBuffer_14_74 : _GEN_3374; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3378 = 4'h1 == lineCounter ? frameBuffer_1_75 : frameBuffer_0_75; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3379 = 4'h2 == lineCounter ? frameBuffer_2_75 : _GEN_3378; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3380 = 4'h3 == lineCounter ? frameBuffer_3_75 : _GEN_3379; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3381 = 4'h4 == lineCounter ? frameBuffer_4_75 : _GEN_3380; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3382 = 4'h5 == lineCounter ? frameBuffer_5_75 : _GEN_3381; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3383 = 4'h6 == lineCounter ? frameBuffer_6_75 : _GEN_3382; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3384 = 4'h7 == lineCounter ? frameBuffer_7_75 : _GEN_3383; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3385 = 4'h8 == lineCounter ? frameBuffer_8_75 : _GEN_3384; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3386 = 4'h9 == lineCounter ? frameBuffer_9_75 : _GEN_3385; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3387 = 4'ha == lineCounter ? frameBuffer_10_75 : _GEN_3386; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3388 = 4'hb == lineCounter ? frameBuffer_11_75 : _GEN_3387; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3389 = 4'hc == lineCounter ? frameBuffer_12_75 : _GEN_3388; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3390 = 4'hd == lineCounter ? frameBuffer_13_75 : _GEN_3389; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3391 = 4'he == lineCounter ? frameBuffer_14_75 : _GEN_3390; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3394 = 4'h1 == lineCounter ? frameBuffer_1_76 : frameBuffer_0_76; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3395 = 4'h2 == lineCounter ? frameBuffer_2_76 : _GEN_3394; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3396 = 4'h3 == lineCounter ? frameBuffer_3_76 : _GEN_3395; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3397 = 4'h4 == lineCounter ? frameBuffer_4_76 : _GEN_3396; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3398 = 4'h5 == lineCounter ? frameBuffer_5_76 : _GEN_3397; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3399 = 4'h6 == lineCounter ? frameBuffer_6_76 : _GEN_3398; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3400 = 4'h7 == lineCounter ? frameBuffer_7_76 : _GEN_3399; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3401 = 4'h8 == lineCounter ? frameBuffer_8_76 : _GEN_3400; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3402 = 4'h9 == lineCounter ? frameBuffer_9_76 : _GEN_3401; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3403 = 4'ha == lineCounter ? frameBuffer_10_76 : _GEN_3402; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3404 = 4'hb == lineCounter ? frameBuffer_11_76 : _GEN_3403; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3405 = 4'hc == lineCounter ? frameBuffer_12_76 : _GEN_3404; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3406 = 4'hd == lineCounter ? frameBuffer_13_76 : _GEN_3405; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3407 = 4'he == lineCounter ? frameBuffer_14_76 : _GEN_3406; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3410 = 4'h1 == lineCounter ? frameBuffer_1_77 : frameBuffer_0_77; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3411 = 4'h2 == lineCounter ? frameBuffer_2_77 : _GEN_3410; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3412 = 4'h3 == lineCounter ? frameBuffer_3_77 : _GEN_3411; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3413 = 4'h4 == lineCounter ? frameBuffer_4_77 : _GEN_3412; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3414 = 4'h5 == lineCounter ? frameBuffer_5_77 : _GEN_3413; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3415 = 4'h6 == lineCounter ? frameBuffer_6_77 : _GEN_3414; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3416 = 4'h7 == lineCounter ? frameBuffer_7_77 : _GEN_3415; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3417 = 4'h8 == lineCounter ? frameBuffer_8_77 : _GEN_3416; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3418 = 4'h9 == lineCounter ? frameBuffer_9_77 : _GEN_3417; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3419 = 4'ha == lineCounter ? frameBuffer_10_77 : _GEN_3418; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3420 = 4'hb == lineCounter ? frameBuffer_11_77 : _GEN_3419; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3421 = 4'hc == lineCounter ? frameBuffer_12_77 : _GEN_3420; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3422 = 4'hd == lineCounter ? frameBuffer_13_77 : _GEN_3421; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3423 = 4'he == lineCounter ? frameBuffer_14_77 : _GEN_3422; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3426 = 4'h1 == lineCounter ? frameBuffer_1_78 : frameBuffer_0_78; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3427 = 4'h2 == lineCounter ? frameBuffer_2_78 : _GEN_3426; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3428 = 4'h3 == lineCounter ? frameBuffer_3_78 : _GEN_3427; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3429 = 4'h4 == lineCounter ? frameBuffer_4_78 : _GEN_3428; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3430 = 4'h5 == lineCounter ? frameBuffer_5_78 : _GEN_3429; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3431 = 4'h6 == lineCounter ? frameBuffer_6_78 : _GEN_3430; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3432 = 4'h7 == lineCounter ? frameBuffer_7_78 : _GEN_3431; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3433 = 4'h8 == lineCounter ? frameBuffer_8_78 : _GEN_3432; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3434 = 4'h9 == lineCounter ? frameBuffer_9_78 : _GEN_3433; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3435 = 4'ha == lineCounter ? frameBuffer_10_78 : _GEN_3434; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3436 = 4'hb == lineCounter ? frameBuffer_11_78 : _GEN_3435; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3437 = 4'hc == lineCounter ? frameBuffer_12_78 : _GEN_3436; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3438 = 4'hd == lineCounter ? frameBuffer_13_78 : _GEN_3437; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3439 = 4'he == lineCounter ? frameBuffer_14_78 : _GEN_3438; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3442 = 4'h1 == lineCounter ? frameBuffer_1_79 : frameBuffer_0_79; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3443 = 4'h2 == lineCounter ? frameBuffer_2_79 : _GEN_3442; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3444 = 4'h3 == lineCounter ? frameBuffer_3_79 : _GEN_3443; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3445 = 4'h4 == lineCounter ? frameBuffer_4_79 : _GEN_3444; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3446 = 4'h5 == lineCounter ? frameBuffer_5_79 : _GEN_3445; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3447 = 4'h6 == lineCounter ? frameBuffer_6_79 : _GEN_3446; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3448 = 4'h7 == lineCounter ? frameBuffer_7_79 : _GEN_3447; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3449 = 4'h8 == lineCounter ? frameBuffer_8_79 : _GEN_3448; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3450 = 4'h9 == lineCounter ? frameBuffer_9_79 : _GEN_3449; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3451 = 4'ha == lineCounter ? frameBuffer_10_79 : _GEN_3450; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3452 = 4'hb == lineCounter ? frameBuffer_11_79 : _GEN_3451; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3453 = 4'hc == lineCounter ? frameBuffer_12_79 : _GEN_3452; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3454 = 4'hd == lineCounter ? frameBuffer_13_79 : _GEN_3453; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3455 = 4'he == lineCounter ? frameBuffer_14_79 : _GEN_3454; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3458 = 4'h1 == lineCounter ? frameBuffer_1_80 : frameBuffer_0_80; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3459 = 4'h2 == lineCounter ? frameBuffer_2_80 : _GEN_3458; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3460 = 4'h3 == lineCounter ? frameBuffer_3_80 : _GEN_3459; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3461 = 4'h4 == lineCounter ? frameBuffer_4_80 : _GEN_3460; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3462 = 4'h5 == lineCounter ? frameBuffer_5_80 : _GEN_3461; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3463 = 4'h6 == lineCounter ? frameBuffer_6_80 : _GEN_3462; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3464 = 4'h7 == lineCounter ? frameBuffer_7_80 : _GEN_3463; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3465 = 4'h8 == lineCounter ? frameBuffer_8_80 : _GEN_3464; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3466 = 4'h9 == lineCounter ? frameBuffer_9_80 : _GEN_3465; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3467 = 4'ha == lineCounter ? frameBuffer_10_80 : _GEN_3466; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3468 = 4'hb == lineCounter ? frameBuffer_11_80 : _GEN_3467; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3469 = 4'hc == lineCounter ? frameBuffer_12_80 : _GEN_3468; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3470 = 4'hd == lineCounter ? frameBuffer_13_80 : _GEN_3469; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3471 = 4'he == lineCounter ? frameBuffer_14_80 : _GEN_3470; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3474 = 4'h1 == lineCounter ? frameBuffer_1_81 : frameBuffer_0_81; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3475 = 4'h2 == lineCounter ? frameBuffer_2_81 : _GEN_3474; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3476 = 4'h3 == lineCounter ? frameBuffer_3_81 : _GEN_3475; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3477 = 4'h4 == lineCounter ? frameBuffer_4_81 : _GEN_3476; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3478 = 4'h5 == lineCounter ? frameBuffer_5_81 : _GEN_3477; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3479 = 4'h6 == lineCounter ? frameBuffer_6_81 : _GEN_3478; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3480 = 4'h7 == lineCounter ? frameBuffer_7_81 : _GEN_3479; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3481 = 4'h8 == lineCounter ? frameBuffer_8_81 : _GEN_3480; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3482 = 4'h9 == lineCounter ? frameBuffer_9_81 : _GEN_3481; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3483 = 4'ha == lineCounter ? frameBuffer_10_81 : _GEN_3482; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3484 = 4'hb == lineCounter ? frameBuffer_11_81 : _GEN_3483; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3485 = 4'hc == lineCounter ? frameBuffer_12_81 : _GEN_3484; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3486 = 4'hd == lineCounter ? frameBuffer_13_81 : _GEN_3485; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3487 = 4'he == lineCounter ? frameBuffer_14_81 : _GEN_3486; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3490 = 4'h1 == lineCounter ? frameBuffer_1_82 : frameBuffer_0_82; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3491 = 4'h2 == lineCounter ? frameBuffer_2_82 : _GEN_3490; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3492 = 4'h3 == lineCounter ? frameBuffer_3_82 : _GEN_3491; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3493 = 4'h4 == lineCounter ? frameBuffer_4_82 : _GEN_3492; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3494 = 4'h5 == lineCounter ? frameBuffer_5_82 : _GEN_3493; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3495 = 4'h6 == lineCounter ? frameBuffer_6_82 : _GEN_3494; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3496 = 4'h7 == lineCounter ? frameBuffer_7_82 : _GEN_3495; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3497 = 4'h8 == lineCounter ? frameBuffer_8_82 : _GEN_3496; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3498 = 4'h9 == lineCounter ? frameBuffer_9_82 : _GEN_3497; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3499 = 4'ha == lineCounter ? frameBuffer_10_82 : _GEN_3498; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3500 = 4'hb == lineCounter ? frameBuffer_11_82 : _GEN_3499; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3501 = 4'hc == lineCounter ? frameBuffer_12_82 : _GEN_3500; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3502 = 4'hd == lineCounter ? frameBuffer_13_82 : _GEN_3501; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3503 = 4'he == lineCounter ? frameBuffer_14_82 : _GEN_3502; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3506 = 4'h1 == lineCounter ? frameBuffer_1_83 : frameBuffer_0_83; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3507 = 4'h2 == lineCounter ? frameBuffer_2_83 : _GEN_3506; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3508 = 4'h3 == lineCounter ? frameBuffer_3_83 : _GEN_3507; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3509 = 4'h4 == lineCounter ? frameBuffer_4_83 : _GEN_3508; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3510 = 4'h5 == lineCounter ? frameBuffer_5_83 : _GEN_3509; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3511 = 4'h6 == lineCounter ? frameBuffer_6_83 : _GEN_3510; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3512 = 4'h7 == lineCounter ? frameBuffer_7_83 : _GEN_3511; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3513 = 4'h8 == lineCounter ? frameBuffer_8_83 : _GEN_3512; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3514 = 4'h9 == lineCounter ? frameBuffer_9_83 : _GEN_3513; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3515 = 4'ha == lineCounter ? frameBuffer_10_83 : _GEN_3514; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3516 = 4'hb == lineCounter ? frameBuffer_11_83 : _GEN_3515; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3517 = 4'hc == lineCounter ? frameBuffer_12_83 : _GEN_3516; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3518 = 4'hd == lineCounter ? frameBuffer_13_83 : _GEN_3517; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3519 = 4'he == lineCounter ? frameBuffer_14_83 : _GEN_3518; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3522 = 4'h1 == lineCounter ? frameBuffer_1_84 : frameBuffer_0_84; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3523 = 4'h2 == lineCounter ? frameBuffer_2_84 : _GEN_3522; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3524 = 4'h3 == lineCounter ? frameBuffer_3_84 : _GEN_3523; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3525 = 4'h4 == lineCounter ? frameBuffer_4_84 : _GEN_3524; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3526 = 4'h5 == lineCounter ? frameBuffer_5_84 : _GEN_3525; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3527 = 4'h6 == lineCounter ? frameBuffer_6_84 : _GEN_3526; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3528 = 4'h7 == lineCounter ? frameBuffer_7_84 : _GEN_3527; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3529 = 4'h8 == lineCounter ? frameBuffer_8_84 : _GEN_3528; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3530 = 4'h9 == lineCounter ? frameBuffer_9_84 : _GEN_3529; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3531 = 4'ha == lineCounter ? frameBuffer_10_84 : _GEN_3530; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3532 = 4'hb == lineCounter ? frameBuffer_11_84 : _GEN_3531; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3533 = 4'hc == lineCounter ? frameBuffer_12_84 : _GEN_3532; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3534 = 4'hd == lineCounter ? frameBuffer_13_84 : _GEN_3533; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3535 = 4'he == lineCounter ? frameBuffer_14_84 : _GEN_3534; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3538 = 4'h1 == lineCounter ? frameBuffer_1_85 : frameBuffer_0_85; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3539 = 4'h2 == lineCounter ? frameBuffer_2_85 : _GEN_3538; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3540 = 4'h3 == lineCounter ? frameBuffer_3_85 : _GEN_3539; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3541 = 4'h4 == lineCounter ? frameBuffer_4_85 : _GEN_3540; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3542 = 4'h5 == lineCounter ? frameBuffer_5_85 : _GEN_3541; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3543 = 4'h6 == lineCounter ? frameBuffer_6_85 : _GEN_3542; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3544 = 4'h7 == lineCounter ? frameBuffer_7_85 : _GEN_3543; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3545 = 4'h8 == lineCounter ? frameBuffer_8_85 : _GEN_3544; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3546 = 4'h9 == lineCounter ? frameBuffer_9_85 : _GEN_3545; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3547 = 4'ha == lineCounter ? frameBuffer_10_85 : _GEN_3546; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3548 = 4'hb == lineCounter ? frameBuffer_11_85 : _GEN_3547; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3549 = 4'hc == lineCounter ? frameBuffer_12_85 : _GEN_3548; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3550 = 4'hd == lineCounter ? frameBuffer_13_85 : _GEN_3549; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3551 = 4'he == lineCounter ? frameBuffer_14_85 : _GEN_3550; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3554 = 4'h1 == lineCounter ? frameBuffer_1_86 : frameBuffer_0_86; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3555 = 4'h2 == lineCounter ? frameBuffer_2_86 : _GEN_3554; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3556 = 4'h3 == lineCounter ? frameBuffer_3_86 : _GEN_3555; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3557 = 4'h4 == lineCounter ? frameBuffer_4_86 : _GEN_3556; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3558 = 4'h5 == lineCounter ? frameBuffer_5_86 : _GEN_3557; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3559 = 4'h6 == lineCounter ? frameBuffer_6_86 : _GEN_3558; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3560 = 4'h7 == lineCounter ? frameBuffer_7_86 : _GEN_3559; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3561 = 4'h8 == lineCounter ? frameBuffer_8_86 : _GEN_3560; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3562 = 4'h9 == lineCounter ? frameBuffer_9_86 : _GEN_3561; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3563 = 4'ha == lineCounter ? frameBuffer_10_86 : _GEN_3562; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3564 = 4'hb == lineCounter ? frameBuffer_11_86 : _GEN_3563; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3565 = 4'hc == lineCounter ? frameBuffer_12_86 : _GEN_3564; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3566 = 4'hd == lineCounter ? frameBuffer_13_86 : _GEN_3565; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3567 = 4'he == lineCounter ? frameBuffer_14_86 : _GEN_3566; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3570 = 4'h1 == lineCounter ? frameBuffer_1_87 : frameBuffer_0_87; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3571 = 4'h2 == lineCounter ? frameBuffer_2_87 : _GEN_3570; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3572 = 4'h3 == lineCounter ? frameBuffer_3_87 : _GEN_3571; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3573 = 4'h4 == lineCounter ? frameBuffer_4_87 : _GEN_3572; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3574 = 4'h5 == lineCounter ? frameBuffer_5_87 : _GEN_3573; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3575 = 4'h6 == lineCounter ? frameBuffer_6_87 : _GEN_3574; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3576 = 4'h7 == lineCounter ? frameBuffer_7_87 : _GEN_3575; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3577 = 4'h8 == lineCounter ? frameBuffer_8_87 : _GEN_3576; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3578 = 4'h9 == lineCounter ? frameBuffer_9_87 : _GEN_3577; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3579 = 4'ha == lineCounter ? frameBuffer_10_87 : _GEN_3578; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3580 = 4'hb == lineCounter ? frameBuffer_11_87 : _GEN_3579; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3581 = 4'hc == lineCounter ? frameBuffer_12_87 : _GEN_3580; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3582 = 4'hd == lineCounter ? frameBuffer_13_87 : _GEN_3581; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3583 = 4'he == lineCounter ? frameBuffer_14_87 : _GEN_3582; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3586 = 4'h1 == lineCounter ? frameBuffer_1_88 : frameBuffer_0_88; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3587 = 4'h2 == lineCounter ? frameBuffer_2_88 : _GEN_3586; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3588 = 4'h3 == lineCounter ? frameBuffer_3_88 : _GEN_3587; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3589 = 4'h4 == lineCounter ? frameBuffer_4_88 : _GEN_3588; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3590 = 4'h5 == lineCounter ? frameBuffer_5_88 : _GEN_3589; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3591 = 4'h6 == lineCounter ? frameBuffer_6_88 : _GEN_3590; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3592 = 4'h7 == lineCounter ? frameBuffer_7_88 : _GEN_3591; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3593 = 4'h8 == lineCounter ? frameBuffer_8_88 : _GEN_3592; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3594 = 4'h9 == lineCounter ? frameBuffer_9_88 : _GEN_3593; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3595 = 4'ha == lineCounter ? frameBuffer_10_88 : _GEN_3594; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3596 = 4'hb == lineCounter ? frameBuffer_11_88 : _GEN_3595; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3597 = 4'hc == lineCounter ? frameBuffer_12_88 : _GEN_3596; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3598 = 4'hd == lineCounter ? frameBuffer_13_88 : _GEN_3597; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3599 = 4'he == lineCounter ? frameBuffer_14_88 : _GEN_3598; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3602 = 4'h1 == lineCounter ? frameBuffer_1_89 : frameBuffer_0_89; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3603 = 4'h2 == lineCounter ? frameBuffer_2_89 : _GEN_3602; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3604 = 4'h3 == lineCounter ? frameBuffer_3_89 : _GEN_3603; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3605 = 4'h4 == lineCounter ? frameBuffer_4_89 : _GEN_3604; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3606 = 4'h5 == lineCounter ? frameBuffer_5_89 : _GEN_3605; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3607 = 4'h6 == lineCounter ? frameBuffer_6_89 : _GEN_3606; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3608 = 4'h7 == lineCounter ? frameBuffer_7_89 : _GEN_3607; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3609 = 4'h8 == lineCounter ? frameBuffer_8_89 : _GEN_3608; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3610 = 4'h9 == lineCounter ? frameBuffer_9_89 : _GEN_3609; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3611 = 4'ha == lineCounter ? frameBuffer_10_89 : _GEN_3610; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3612 = 4'hb == lineCounter ? frameBuffer_11_89 : _GEN_3611; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3613 = 4'hc == lineCounter ? frameBuffer_12_89 : _GEN_3612; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3614 = 4'hd == lineCounter ? frameBuffer_13_89 : _GEN_3613; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3615 = 4'he == lineCounter ? frameBuffer_14_89 : _GEN_3614; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3618 = 4'h1 == lineCounter ? frameBuffer_1_90 : frameBuffer_0_90; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3619 = 4'h2 == lineCounter ? frameBuffer_2_90 : _GEN_3618; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3620 = 4'h3 == lineCounter ? frameBuffer_3_90 : _GEN_3619; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3621 = 4'h4 == lineCounter ? frameBuffer_4_90 : _GEN_3620; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3622 = 4'h5 == lineCounter ? frameBuffer_5_90 : _GEN_3621; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3623 = 4'h6 == lineCounter ? frameBuffer_6_90 : _GEN_3622; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3624 = 4'h7 == lineCounter ? frameBuffer_7_90 : _GEN_3623; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3625 = 4'h8 == lineCounter ? frameBuffer_8_90 : _GEN_3624; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3626 = 4'h9 == lineCounter ? frameBuffer_9_90 : _GEN_3625; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3627 = 4'ha == lineCounter ? frameBuffer_10_90 : _GEN_3626; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3628 = 4'hb == lineCounter ? frameBuffer_11_90 : _GEN_3627; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3629 = 4'hc == lineCounter ? frameBuffer_12_90 : _GEN_3628; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3630 = 4'hd == lineCounter ? frameBuffer_13_90 : _GEN_3629; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3631 = 4'he == lineCounter ? frameBuffer_14_90 : _GEN_3630; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3634 = 4'h1 == lineCounter ? frameBuffer_1_91 : frameBuffer_0_91; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3635 = 4'h2 == lineCounter ? frameBuffer_2_91 : _GEN_3634; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3636 = 4'h3 == lineCounter ? frameBuffer_3_91 : _GEN_3635; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3637 = 4'h4 == lineCounter ? frameBuffer_4_91 : _GEN_3636; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3638 = 4'h5 == lineCounter ? frameBuffer_5_91 : _GEN_3637; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3639 = 4'h6 == lineCounter ? frameBuffer_6_91 : _GEN_3638; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3640 = 4'h7 == lineCounter ? frameBuffer_7_91 : _GEN_3639; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3641 = 4'h8 == lineCounter ? frameBuffer_8_91 : _GEN_3640; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3642 = 4'h9 == lineCounter ? frameBuffer_9_91 : _GEN_3641; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3643 = 4'ha == lineCounter ? frameBuffer_10_91 : _GEN_3642; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3644 = 4'hb == lineCounter ? frameBuffer_11_91 : _GEN_3643; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3645 = 4'hc == lineCounter ? frameBuffer_12_91 : _GEN_3644; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3646 = 4'hd == lineCounter ? frameBuffer_13_91 : _GEN_3645; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3647 = 4'he == lineCounter ? frameBuffer_14_91 : _GEN_3646; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3650 = 4'h1 == lineCounter ? frameBuffer_1_92 : frameBuffer_0_92; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3651 = 4'h2 == lineCounter ? frameBuffer_2_92 : _GEN_3650; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3652 = 4'h3 == lineCounter ? frameBuffer_3_92 : _GEN_3651; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3653 = 4'h4 == lineCounter ? frameBuffer_4_92 : _GEN_3652; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3654 = 4'h5 == lineCounter ? frameBuffer_5_92 : _GEN_3653; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3655 = 4'h6 == lineCounter ? frameBuffer_6_92 : _GEN_3654; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3656 = 4'h7 == lineCounter ? frameBuffer_7_92 : _GEN_3655; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3657 = 4'h8 == lineCounter ? frameBuffer_8_92 : _GEN_3656; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3658 = 4'h9 == lineCounter ? frameBuffer_9_92 : _GEN_3657; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3659 = 4'ha == lineCounter ? frameBuffer_10_92 : _GEN_3658; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3660 = 4'hb == lineCounter ? frameBuffer_11_92 : _GEN_3659; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3661 = 4'hc == lineCounter ? frameBuffer_12_92 : _GEN_3660; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3662 = 4'hd == lineCounter ? frameBuffer_13_92 : _GEN_3661; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3663 = 4'he == lineCounter ? frameBuffer_14_92 : _GEN_3662; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3666 = 4'h1 == lineCounter ? frameBuffer_1_93 : frameBuffer_0_93; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3667 = 4'h2 == lineCounter ? frameBuffer_2_93 : _GEN_3666; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3668 = 4'h3 == lineCounter ? frameBuffer_3_93 : _GEN_3667; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3669 = 4'h4 == lineCounter ? frameBuffer_4_93 : _GEN_3668; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3670 = 4'h5 == lineCounter ? frameBuffer_5_93 : _GEN_3669; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3671 = 4'h6 == lineCounter ? frameBuffer_6_93 : _GEN_3670; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3672 = 4'h7 == lineCounter ? frameBuffer_7_93 : _GEN_3671; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3673 = 4'h8 == lineCounter ? frameBuffer_8_93 : _GEN_3672; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3674 = 4'h9 == lineCounter ? frameBuffer_9_93 : _GEN_3673; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3675 = 4'ha == lineCounter ? frameBuffer_10_93 : _GEN_3674; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3676 = 4'hb == lineCounter ? frameBuffer_11_93 : _GEN_3675; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3677 = 4'hc == lineCounter ? frameBuffer_12_93 : _GEN_3676; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3678 = 4'hd == lineCounter ? frameBuffer_13_93 : _GEN_3677; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3679 = 4'he == lineCounter ? frameBuffer_14_93 : _GEN_3678; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3682 = 4'h1 == lineCounter ? frameBuffer_1_94 : frameBuffer_0_94; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3683 = 4'h2 == lineCounter ? frameBuffer_2_94 : _GEN_3682; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3684 = 4'h3 == lineCounter ? frameBuffer_3_94 : _GEN_3683; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3685 = 4'h4 == lineCounter ? frameBuffer_4_94 : _GEN_3684; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3686 = 4'h5 == lineCounter ? frameBuffer_5_94 : _GEN_3685; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3687 = 4'h6 == lineCounter ? frameBuffer_6_94 : _GEN_3686; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3688 = 4'h7 == lineCounter ? frameBuffer_7_94 : _GEN_3687; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3689 = 4'h8 == lineCounter ? frameBuffer_8_94 : _GEN_3688; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3690 = 4'h9 == lineCounter ? frameBuffer_9_94 : _GEN_3689; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3691 = 4'ha == lineCounter ? frameBuffer_10_94 : _GEN_3690; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3692 = 4'hb == lineCounter ? frameBuffer_11_94 : _GEN_3691; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3693 = 4'hc == lineCounter ? frameBuffer_12_94 : _GEN_3692; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3694 = 4'hd == lineCounter ? frameBuffer_13_94 : _GEN_3693; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3695 = 4'he == lineCounter ? frameBuffer_14_94 : _GEN_3694; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3698 = 4'h1 == lineCounter ? frameBuffer_1_95 : frameBuffer_0_95; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3699 = 4'h2 == lineCounter ? frameBuffer_2_95 : _GEN_3698; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3700 = 4'h3 == lineCounter ? frameBuffer_3_95 : _GEN_3699; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3701 = 4'h4 == lineCounter ? frameBuffer_4_95 : _GEN_3700; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3702 = 4'h5 == lineCounter ? frameBuffer_5_95 : _GEN_3701; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3703 = 4'h6 == lineCounter ? frameBuffer_6_95 : _GEN_3702; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3704 = 4'h7 == lineCounter ? frameBuffer_7_95 : _GEN_3703; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3705 = 4'h8 == lineCounter ? frameBuffer_8_95 : _GEN_3704; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3706 = 4'h9 == lineCounter ? frameBuffer_9_95 : _GEN_3705; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3707 = 4'ha == lineCounter ? frameBuffer_10_95 : _GEN_3706; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3708 = 4'hb == lineCounter ? frameBuffer_11_95 : _GEN_3707; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3709 = 4'hc == lineCounter ? frameBuffer_12_95 : _GEN_3708; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3710 = 4'hd == lineCounter ? frameBuffer_13_95 : _GEN_3709; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3711 = 4'he == lineCounter ? frameBuffer_14_95 : _GEN_3710; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3714 = 4'h1 == lineCounter ? frameBuffer_1_96 : frameBuffer_0_96; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3715 = 4'h2 == lineCounter ? frameBuffer_2_96 : _GEN_3714; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3716 = 4'h3 == lineCounter ? frameBuffer_3_96 : _GEN_3715; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3717 = 4'h4 == lineCounter ? frameBuffer_4_96 : _GEN_3716; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3718 = 4'h5 == lineCounter ? frameBuffer_5_96 : _GEN_3717; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3719 = 4'h6 == lineCounter ? frameBuffer_6_96 : _GEN_3718; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3720 = 4'h7 == lineCounter ? frameBuffer_7_96 : _GEN_3719; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3721 = 4'h8 == lineCounter ? frameBuffer_8_96 : _GEN_3720; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3722 = 4'h9 == lineCounter ? frameBuffer_9_96 : _GEN_3721; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3723 = 4'ha == lineCounter ? frameBuffer_10_96 : _GEN_3722; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3724 = 4'hb == lineCounter ? frameBuffer_11_96 : _GEN_3723; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3725 = 4'hc == lineCounter ? frameBuffer_12_96 : _GEN_3724; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3726 = 4'hd == lineCounter ? frameBuffer_13_96 : _GEN_3725; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3727 = 4'he == lineCounter ? frameBuffer_14_96 : _GEN_3726; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3730 = 4'h1 == lineCounter ? frameBuffer_1_97 : frameBuffer_0_97; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3731 = 4'h2 == lineCounter ? frameBuffer_2_97 : _GEN_3730; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3732 = 4'h3 == lineCounter ? frameBuffer_3_97 : _GEN_3731; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3733 = 4'h4 == lineCounter ? frameBuffer_4_97 : _GEN_3732; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3734 = 4'h5 == lineCounter ? frameBuffer_5_97 : _GEN_3733; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3735 = 4'h6 == lineCounter ? frameBuffer_6_97 : _GEN_3734; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3736 = 4'h7 == lineCounter ? frameBuffer_7_97 : _GEN_3735; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3737 = 4'h8 == lineCounter ? frameBuffer_8_97 : _GEN_3736; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3738 = 4'h9 == lineCounter ? frameBuffer_9_97 : _GEN_3737; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3739 = 4'ha == lineCounter ? frameBuffer_10_97 : _GEN_3738; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3740 = 4'hb == lineCounter ? frameBuffer_11_97 : _GEN_3739; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3741 = 4'hc == lineCounter ? frameBuffer_12_97 : _GEN_3740; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3742 = 4'hd == lineCounter ? frameBuffer_13_97 : _GEN_3741; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3743 = 4'he == lineCounter ? frameBuffer_14_97 : _GEN_3742; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3746 = 4'h1 == lineCounter ? frameBuffer_1_98 : frameBuffer_0_98; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3747 = 4'h2 == lineCounter ? frameBuffer_2_98 : _GEN_3746; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3748 = 4'h3 == lineCounter ? frameBuffer_3_98 : _GEN_3747; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3749 = 4'h4 == lineCounter ? frameBuffer_4_98 : _GEN_3748; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3750 = 4'h5 == lineCounter ? frameBuffer_5_98 : _GEN_3749; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3751 = 4'h6 == lineCounter ? frameBuffer_6_98 : _GEN_3750; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3752 = 4'h7 == lineCounter ? frameBuffer_7_98 : _GEN_3751; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3753 = 4'h8 == lineCounter ? frameBuffer_8_98 : _GEN_3752; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3754 = 4'h9 == lineCounter ? frameBuffer_9_98 : _GEN_3753; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3755 = 4'ha == lineCounter ? frameBuffer_10_98 : _GEN_3754; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3756 = 4'hb == lineCounter ? frameBuffer_11_98 : _GEN_3755; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3757 = 4'hc == lineCounter ? frameBuffer_12_98 : _GEN_3756; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3758 = 4'hd == lineCounter ? frameBuffer_13_98 : _GEN_3757; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3759 = 4'he == lineCounter ? frameBuffer_14_98 : _GEN_3758; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3762 = 4'h1 == lineCounter ? frameBuffer_1_99 : frameBuffer_0_99; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3763 = 4'h2 == lineCounter ? frameBuffer_2_99 : _GEN_3762; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3764 = 4'h3 == lineCounter ? frameBuffer_3_99 : _GEN_3763; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3765 = 4'h4 == lineCounter ? frameBuffer_4_99 : _GEN_3764; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3766 = 4'h5 == lineCounter ? frameBuffer_5_99 : _GEN_3765; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3767 = 4'h6 == lineCounter ? frameBuffer_6_99 : _GEN_3766; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3768 = 4'h7 == lineCounter ? frameBuffer_7_99 : _GEN_3767; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3769 = 4'h8 == lineCounter ? frameBuffer_8_99 : _GEN_3768; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3770 = 4'h9 == lineCounter ? frameBuffer_9_99 : _GEN_3769; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3771 = 4'ha == lineCounter ? frameBuffer_10_99 : _GEN_3770; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3772 = 4'hb == lineCounter ? frameBuffer_11_99 : _GEN_3771; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3773 = 4'hc == lineCounter ? frameBuffer_12_99 : _GEN_3772; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3774 = 4'hd == lineCounter ? frameBuffer_13_99 : _GEN_3773; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3775 = 4'he == lineCounter ? frameBuffer_14_99 : _GEN_3774; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3778 = 4'h1 == lineCounter ? frameBuffer_1_100 : frameBuffer_0_100; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3779 = 4'h2 == lineCounter ? frameBuffer_2_100 : _GEN_3778; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3780 = 4'h3 == lineCounter ? frameBuffer_3_100 : _GEN_3779; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3781 = 4'h4 == lineCounter ? frameBuffer_4_100 : _GEN_3780; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3782 = 4'h5 == lineCounter ? frameBuffer_5_100 : _GEN_3781; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3783 = 4'h6 == lineCounter ? frameBuffer_6_100 : _GEN_3782; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3784 = 4'h7 == lineCounter ? frameBuffer_7_100 : _GEN_3783; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3785 = 4'h8 == lineCounter ? frameBuffer_8_100 : _GEN_3784; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3786 = 4'h9 == lineCounter ? frameBuffer_9_100 : _GEN_3785; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3787 = 4'ha == lineCounter ? frameBuffer_10_100 : _GEN_3786; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3788 = 4'hb == lineCounter ? frameBuffer_11_100 : _GEN_3787; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3789 = 4'hc == lineCounter ? frameBuffer_12_100 : _GEN_3788; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3790 = 4'hd == lineCounter ? frameBuffer_13_100 : _GEN_3789; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3791 = 4'he == lineCounter ? frameBuffer_14_100 : _GEN_3790; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3794 = 4'h1 == lineCounter ? frameBuffer_1_101 : frameBuffer_0_101; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3795 = 4'h2 == lineCounter ? frameBuffer_2_101 : _GEN_3794; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3796 = 4'h3 == lineCounter ? frameBuffer_3_101 : _GEN_3795; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3797 = 4'h4 == lineCounter ? frameBuffer_4_101 : _GEN_3796; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3798 = 4'h5 == lineCounter ? frameBuffer_5_101 : _GEN_3797; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3799 = 4'h6 == lineCounter ? frameBuffer_6_101 : _GEN_3798; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3800 = 4'h7 == lineCounter ? frameBuffer_7_101 : _GEN_3799; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3801 = 4'h8 == lineCounter ? frameBuffer_8_101 : _GEN_3800; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3802 = 4'h9 == lineCounter ? frameBuffer_9_101 : _GEN_3801; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3803 = 4'ha == lineCounter ? frameBuffer_10_101 : _GEN_3802; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3804 = 4'hb == lineCounter ? frameBuffer_11_101 : _GEN_3803; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3805 = 4'hc == lineCounter ? frameBuffer_12_101 : _GEN_3804; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3806 = 4'hd == lineCounter ? frameBuffer_13_101 : _GEN_3805; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3807 = 4'he == lineCounter ? frameBuffer_14_101 : _GEN_3806; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3810 = 4'h1 == lineCounter ? frameBuffer_1_102 : frameBuffer_0_102; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3811 = 4'h2 == lineCounter ? frameBuffer_2_102 : _GEN_3810; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3812 = 4'h3 == lineCounter ? frameBuffer_3_102 : _GEN_3811; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3813 = 4'h4 == lineCounter ? frameBuffer_4_102 : _GEN_3812; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3814 = 4'h5 == lineCounter ? frameBuffer_5_102 : _GEN_3813; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3815 = 4'h6 == lineCounter ? frameBuffer_6_102 : _GEN_3814; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3816 = 4'h7 == lineCounter ? frameBuffer_7_102 : _GEN_3815; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3817 = 4'h8 == lineCounter ? frameBuffer_8_102 : _GEN_3816; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3818 = 4'h9 == lineCounter ? frameBuffer_9_102 : _GEN_3817; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3819 = 4'ha == lineCounter ? frameBuffer_10_102 : _GEN_3818; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3820 = 4'hb == lineCounter ? frameBuffer_11_102 : _GEN_3819; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3821 = 4'hc == lineCounter ? frameBuffer_12_102 : _GEN_3820; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3822 = 4'hd == lineCounter ? frameBuffer_13_102 : _GEN_3821; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3823 = 4'he == lineCounter ? frameBuffer_14_102 : _GEN_3822; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3826 = 4'h1 == lineCounter ? frameBuffer_1_103 : frameBuffer_0_103; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3827 = 4'h2 == lineCounter ? frameBuffer_2_103 : _GEN_3826; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3828 = 4'h3 == lineCounter ? frameBuffer_3_103 : _GEN_3827; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3829 = 4'h4 == lineCounter ? frameBuffer_4_103 : _GEN_3828; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3830 = 4'h5 == lineCounter ? frameBuffer_5_103 : _GEN_3829; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3831 = 4'h6 == lineCounter ? frameBuffer_6_103 : _GEN_3830; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3832 = 4'h7 == lineCounter ? frameBuffer_7_103 : _GEN_3831; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3833 = 4'h8 == lineCounter ? frameBuffer_8_103 : _GEN_3832; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3834 = 4'h9 == lineCounter ? frameBuffer_9_103 : _GEN_3833; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3835 = 4'ha == lineCounter ? frameBuffer_10_103 : _GEN_3834; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3836 = 4'hb == lineCounter ? frameBuffer_11_103 : _GEN_3835; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3837 = 4'hc == lineCounter ? frameBuffer_12_103 : _GEN_3836; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3838 = 4'hd == lineCounter ? frameBuffer_13_103 : _GEN_3837; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3839 = 4'he == lineCounter ? frameBuffer_14_103 : _GEN_3838; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3842 = 4'h1 == lineCounter ? frameBuffer_1_104 : frameBuffer_0_104; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3843 = 4'h2 == lineCounter ? frameBuffer_2_104 : _GEN_3842; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3844 = 4'h3 == lineCounter ? frameBuffer_3_104 : _GEN_3843; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3845 = 4'h4 == lineCounter ? frameBuffer_4_104 : _GEN_3844; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3846 = 4'h5 == lineCounter ? frameBuffer_5_104 : _GEN_3845; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3847 = 4'h6 == lineCounter ? frameBuffer_6_104 : _GEN_3846; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3848 = 4'h7 == lineCounter ? frameBuffer_7_104 : _GEN_3847; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3849 = 4'h8 == lineCounter ? frameBuffer_8_104 : _GEN_3848; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3850 = 4'h9 == lineCounter ? frameBuffer_9_104 : _GEN_3849; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3851 = 4'ha == lineCounter ? frameBuffer_10_104 : _GEN_3850; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3852 = 4'hb == lineCounter ? frameBuffer_11_104 : _GEN_3851; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3853 = 4'hc == lineCounter ? frameBuffer_12_104 : _GEN_3852; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3854 = 4'hd == lineCounter ? frameBuffer_13_104 : _GEN_3853; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3855 = 4'he == lineCounter ? frameBuffer_14_104 : _GEN_3854; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3858 = 4'h1 == lineCounter ? frameBuffer_1_105 : frameBuffer_0_105; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3859 = 4'h2 == lineCounter ? frameBuffer_2_105 : _GEN_3858; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3860 = 4'h3 == lineCounter ? frameBuffer_3_105 : _GEN_3859; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3861 = 4'h4 == lineCounter ? frameBuffer_4_105 : _GEN_3860; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3862 = 4'h5 == lineCounter ? frameBuffer_5_105 : _GEN_3861; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3863 = 4'h6 == lineCounter ? frameBuffer_6_105 : _GEN_3862; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3864 = 4'h7 == lineCounter ? frameBuffer_7_105 : _GEN_3863; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3865 = 4'h8 == lineCounter ? frameBuffer_8_105 : _GEN_3864; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3866 = 4'h9 == lineCounter ? frameBuffer_9_105 : _GEN_3865; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3867 = 4'ha == lineCounter ? frameBuffer_10_105 : _GEN_3866; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3868 = 4'hb == lineCounter ? frameBuffer_11_105 : _GEN_3867; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3869 = 4'hc == lineCounter ? frameBuffer_12_105 : _GEN_3868; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3870 = 4'hd == lineCounter ? frameBuffer_13_105 : _GEN_3869; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3871 = 4'he == lineCounter ? frameBuffer_14_105 : _GEN_3870; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3874 = 4'h1 == lineCounter ? frameBuffer_1_106 : frameBuffer_0_106; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3875 = 4'h2 == lineCounter ? frameBuffer_2_106 : _GEN_3874; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3876 = 4'h3 == lineCounter ? frameBuffer_3_106 : _GEN_3875; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3877 = 4'h4 == lineCounter ? frameBuffer_4_106 : _GEN_3876; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3878 = 4'h5 == lineCounter ? frameBuffer_5_106 : _GEN_3877; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3879 = 4'h6 == lineCounter ? frameBuffer_6_106 : _GEN_3878; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3880 = 4'h7 == lineCounter ? frameBuffer_7_106 : _GEN_3879; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3881 = 4'h8 == lineCounter ? frameBuffer_8_106 : _GEN_3880; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3882 = 4'h9 == lineCounter ? frameBuffer_9_106 : _GEN_3881; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3883 = 4'ha == lineCounter ? frameBuffer_10_106 : _GEN_3882; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3884 = 4'hb == lineCounter ? frameBuffer_11_106 : _GEN_3883; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3885 = 4'hc == lineCounter ? frameBuffer_12_106 : _GEN_3884; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3886 = 4'hd == lineCounter ? frameBuffer_13_106 : _GEN_3885; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3887 = 4'he == lineCounter ? frameBuffer_14_106 : _GEN_3886; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3890 = 4'h1 == lineCounter ? frameBuffer_1_107 : frameBuffer_0_107; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3891 = 4'h2 == lineCounter ? frameBuffer_2_107 : _GEN_3890; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3892 = 4'h3 == lineCounter ? frameBuffer_3_107 : _GEN_3891; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3893 = 4'h4 == lineCounter ? frameBuffer_4_107 : _GEN_3892; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3894 = 4'h5 == lineCounter ? frameBuffer_5_107 : _GEN_3893; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3895 = 4'h6 == lineCounter ? frameBuffer_6_107 : _GEN_3894; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3896 = 4'h7 == lineCounter ? frameBuffer_7_107 : _GEN_3895; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3897 = 4'h8 == lineCounter ? frameBuffer_8_107 : _GEN_3896; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3898 = 4'h9 == lineCounter ? frameBuffer_9_107 : _GEN_3897; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3899 = 4'ha == lineCounter ? frameBuffer_10_107 : _GEN_3898; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3900 = 4'hb == lineCounter ? frameBuffer_11_107 : _GEN_3899; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3901 = 4'hc == lineCounter ? frameBuffer_12_107 : _GEN_3900; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3902 = 4'hd == lineCounter ? frameBuffer_13_107 : _GEN_3901; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3903 = 4'he == lineCounter ? frameBuffer_14_107 : _GEN_3902; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3906 = 4'h1 == lineCounter ? frameBuffer_1_108 : frameBuffer_0_108; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3907 = 4'h2 == lineCounter ? frameBuffer_2_108 : _GEN_3906; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3908 = 4'h3 == lineCounter ? frameBuffer_3_108 : _GEN_3907; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3909 = 4'h4 == lineCounter ? frameBuffer_4_108 : _GEN_3908; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3910 = 4'h5 == lineCounter ? frameBuffer_5_108 : _GEN_3909; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3911 = 4'h6 == lineCounter ? frameBuffer_6_108 : _GEN_3910; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3912 = 4'h7 == lineCounter ? frameBuffer_7_108 : _GEN_3911; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3913 = 4'h8 == lineCounter ? frameBuffer_8_108 : _GEN_3912; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3914 = 4'h9 == lineCounter ? frameBuffer_9_108 : _GEN_3913; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3915 = 4'ha == lineCounter ? frameBuffer_10_108 : _GEN_3914; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3916 = 4'hb == lineCounter ? frameBuffer_11_108 : _GEN_3915; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3917 = 4'hc == lineCounter ? frameBuffer_12_108 : _GEN_3916; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3918 = 4'hd == lineCounter ? frameBuffer_13_108 : _GEN_3917; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3919 = 4'he == lineCounter ? frameBuffer_14_108 : _GEN_3918; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3922 = 4'h1 == lineCounter ? frameBuffer_1_109 : frameBuffer_0_109; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3923 = 4'h2 == lineCounter ? frameBuffer_2_109 : _GEN_3922; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3924 = 4'h3 == lineCounter ? frameBuffer_3_109 : _GEN_3923; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3925 = 4'h4 == lineCounter ? frameBuffer_4_109 : _GEN_3924; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3926 = 4'h5 == lineCounter ? frameBuffer_5_109 : _GEN_3925; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3927 = 4'h6 == lineCounter ? frameBuffer_6_109 : _GEN_3926; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3928 = 4'h7 == lineCounter ? frameBuffer_7_109 : _GEN_3927; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3929 = 4'h8 == lineCounter ? frameBuffer_8_109 : _GEN_3928; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3930 = 4'h9 == lineCounter ? frameBuffer_9_109 : _GEN_3929; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3931 = 4'ha == lineCounter ? frameBuffer_10_109 : _GEN_3930; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3932 = 4'hb == lineCounter ? frameBuffer_11_109 : _GEN_3931; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3933 = 4'hc == lineCounter ? frameBuffer_12_109 : _GEN_3932; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3934 = 4'hd == lineCounter ? frameBuffer_13_109 : _GEN_3933; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3935 = 4'he == lineCounter ? frameBuffer_14_109 : _GEN_3934; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3938 = 4'h1 == lineCounter ? frameBuffer_1_110 : frameBuffer_0_110; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3939 = 4'h2 == lineCounter ? frameBuffer_2_110 : _GEN_3938; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3940 = 4'h3 == lineCounter ? frameBuffer_3_110 : _GEN_3939; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3941 = 4'h4 == lineCounter ? frameBuffer_4_110 : _GEN_3940; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3942 = 4'h5 == lineCounter ? frameBuffer_5_110 : _GEN_3941; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3943 = 4'h6 == lineCounter ? frameBuffer_6_110 : _GEN_3942; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3944 = 4'h7 == lineCounter ? frameBuffer_7_110 : _GEN_3943; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3945 = 4'h8 == lineCounter ? frameBuffer_8_110 : _GEN_3944; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3946 = 4'h9 == lineCounter ? frameBuffer_9_110 : _GEN_3945; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3947 = 4'ha == lineCounter ? frameBuffer_10_110 : _GEN_3946; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3948 = 4'hb == lineCounter ? frameBuffer_11_110 : _GEN_3947; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3949 = 4'hc == lineCounter ? frameBuffer_12_110 : _GEN_3948; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3950 = 4'hd == lineCounter ? frameBuffer_13_110 : _GEN_3949; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3951 = 4'he == lineCounter ? frameBuffer_14_110 : _GEN_3950; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3954 = 4'h1 == lineCounter ? frameBuffer_1_111 : frameBuffer_0_111; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3955 = 4'h2 == lineCounter ? frameBuffer_2_111 : _GEN_3954; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3956 = 4'h3 == lineCounter ? frameBuffer_3_111 : _GEN_3955; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3957 = 4'h4 == lineCounter ? frameBuffer_4_111 : _GEN_3956; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3958 = 4'h5 == lineCounter ? frameBuffer_5_111 : _GEN_3957; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3959 = 4'h6 == lineCounter ? frameBuffer_6_111 : _GEN_3958; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3960 = 4'h7 == lineCounter ? frameBuffer_7_111 : _GEN_3959; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3961 = 4'h8 == lineCounter ? frameBuffer_8_111 : _GEN_3960; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3962 = 4'h9 == lineCounter ? frameBuffer_9_111 : _GEN_3961; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3963 = 4'ha == lineCounter ? frameBuffer_10_111 : _GEN_3962; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3964 = 4'hb == lineCounter ? frameBuffer_11_111 : _GEN_3963; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3965 = 4'hc == lineCounter ? frameBuffer_12_111 : _GEN_3964; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3966 = 4'hd == lineCounter ? frameBuffer_13_111 : _GEN_3965; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3967 = 4'he == lineCounter ? frameBuffer_14_111 : _GEN_3966; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3970 = 4'h1 == lineCounter ? frameBuffer_1_112 : frameBuffer_0_112; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3971 = 4'h2 == lineCounter ? frameBuffer_2_112 : _GEN_3970; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3972 = 4'h3 == lineCounter ? frameBuffer_3_112 : _GEN_3971; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3973 = 4'h4 == lineCounter ? frameBuffer_4_112 : _GEN_3972; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3974 = 4'h5 == lineCounter ? frameBuffer_5_112 : _GEN_3973; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3975 = 4'h6 == lineCounter ? frameBuffer_6_112 : _GEN_3974; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3976 = 4'h7 == lineCounter ? frameBuffer_7_112 : _GEN_3975; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3977 = 4'h8 == lineCounter ? frameBuffer_8_112 : _GEN_3976; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3978 = 4'h9 == lineCounter ? frameBuffer_9_112 : _GEN_3977; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3979 = 4'ha == lineCounter ? frameBuffer_10_112 : _GEN_3978; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3980 = 4'hb == lineCounter ? frameBuffer_11_112 : _GEN_3979; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3981 = 4'hc == lineCounter ? frameBuffer_12_112 : _GEN_3980; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3982 = 4'hd == lineCounter ? frameBuffer_13_112 : _GEN_3981; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3983 = 4'he == lineCounter ? frameBuffer_14_112 : _GEN_3982; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3986 = 4'h1 == lineCounter ? frameBuffer_1_113 : frameBuffer_0_113; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3987 = 4'h2 == lineCounter ? frameBuffer_2_113 : _GEN_3986; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3988 = 4'h3 == lineCounter ? frameBuffer_3_113 : _GEN_3987; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3989 = 4'h4 == lineCounter ? frameBuffer_4_113 : _GEN_3988; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3990 = 4'h5 == lineCounter ? frameBuffer_5_113 : _GEN_3989; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3991 = 4'h6 == lineCounter ? frameBuffer_6_113 : _GEN_3990; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3992 = 4'h7 == lineCounter ? frameBuffer_7_113 : _GEN_3991; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3993 = 4'h8 == lineCounter ? frameBuffer_8_113 : _GEN_3992; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3994 = 4'h9 == lineCounter ? frameBuffer_9_113 : _GEN_3993; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3995 = 4'ha == lineCounter ? frameBuffer_10_113 : _GEN_3994; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3996 = 4'hb == lineCounter ? frameBuffer_11_113 : _GEN_3995; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3997 = 4'hc == lineCounter ? frameBuffer_12_113 : _GEN_3996; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3998 = 4'hd == lineCounter ? frameBuffer_13_113 : _GEN_3997; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_3999 = 4'he == lineCounter ? frameBuffer_14_113 : _GEN_3998; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4002 = 4'h1 == lineCounter ? frameBuffer_1_114 : frameBuffer_0_114; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4003 = 4'h2 == lineCounter ? frameBuffer_2_114 : _GEN_4002; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4004 = 4'h3 == lineCounter ? frameBuffer_3_114 : _GEN_4003; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4005 = 4'h4 == lineCounter ? frameBuffer_4_114 : _GEN_4004; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4006 = 4'h5 == lineCounter ? frameBuffer_5_114 : _GEN_4005; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4007 = 4'h6 == lineCounter ? frameBuffer_6_114 : _GEN_4006; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4008 = 4'h7 == lineCounter ? frameBuffer_7_114 : _GEN_4007; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4009 = 4'h8 == lineCounter ? frameBuffer_8_114 : _GEN_4008; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4010 = 4'h9 == lineCounter ? frameBuffer_9_114 : _GEN_4009; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4011 = 4'ha == lineCounter ? frameBuffer_10_114 : _GEN_4010; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4012 = 4'hb == lineCounter ? frameBuffer_11_114 : _GEN_4011; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4013 = 4'hc == lineCounter ? frameBuffer_12_114 : _GEN_4012; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4014 = 4'hd == lineCounter ? frameBuffer_13_114 : _GEN_4013; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4015 = 4'he == lineCounter ? frameBuffer_14_114 : _GEN_4014; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4018 = 4'h1 == lineCounter ? frameBuffer_1_115 : frameBuffer_0_115; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4019 = 4'h2 == lineCounter ? frameBuffer_2_115 : _GEN_4018; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4020 = 4'h3 == lineCounter ? frameBuffer_3_115 : _GEN_4019; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4021 = 4'h4 == lineCounter ? frameBuffer_4_115 : _GEN_4020; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4022 = 4'h5 == lineCounter ? frameBuffer_5_115 : _GEN_4021; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4023 = 4'h6 == lineCounter ? frameBuffer_6_115 : _GEN_4022; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4024 = 4'h7 == lineCounter ? frameBuffer_7_115 : _GEN_4023; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4025 = 4'h8 == lineCounter ? frameBuffer_8_115 : _GEN_4024; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4026 = 4'h9 == lineCounter ? frameBuffer_9_115 : _GEN_4025; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4027 = 4'ha == lineCounter ? frameBuffer_10_115 : _GEN_4026; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4028 = 4'hb == lineCounter ? frameBuffer_11_115 : _GEN_4027; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4029 = 4'hc == lineCounter ? frameBuffer_12_115 : _GEN_4028; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4030 = 4'hd == lineCounter ? frameBuffer_13_115 : _GEN_4029; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4031 = 4'he == lineCounter ? frameBuffer_14_115 : _GEN_4030; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4034 = 4'h1 == lineCounter ? frameBuffer_1_116 : frameBuffer_0_116; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4035 = 4'h2 == lineCounter ? frameBuffer_2_116 : _GEN_4034; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4036 = 4'h3 == lineCounter ? frameBuffer_3_116 : _GEN_4035; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4037 = 4'h4 == lineCounter ? frameBuffer_4_116 : _GEN_4036; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4038 = 4'h5 == lineCounter ? frameBuffer_5_116 : _GEN_4037; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4039 = 4'h6 == lineCounter ? frameBuffer_6_116 : _GEN_4038; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4040 = 4'h7 == lineCounter ? frameBuffer_7_116 : _GEN_4039; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4041 = 4'h8 == lineCounter ? frameBuffer_8_116 : _GEN_4040; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4042 = 4'h9 == lineCounter ? frameBuffer_9_116 : _GEN_4041; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4043 = 4'ha == lineCounter ? frameBuffer_10_116 : _GEN_4042; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4044 = 4'hb == lineCounter ? frameBuffer_11_116 : _GEN_4043; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4045 = 4'hc == lineCounter ? frameBuffer_12_116 : _GEN_4044; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4046 = 4'hd == lineCounter ? frameBuffer_13_116 : _GEN_4045; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4047 = 4'he == lineCounter ? frameBuffer_14_116 : _GEN_4046; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4050 = 4'h1 == lineCounter ? frameBuffer_1_117 : frameBuffer_0_117; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4051 = 4'h2 == lineCounter ? frameBuffer_2_117 : _GEN_4050; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4052 = 4'h3 == lineCounter ? frameBuffer_3_117 : _GEN_4051; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4053 = 4'h4 == lineCounter ? frameBuffer_4_117 : _GEN_4052; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4054 = 4'h5 == lineCounter ? frameBuffer_5_117 : _GEN_4053; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4055 = 4'h6 == lineCounter ? frameBuffer_6_117 : _GEN_4054; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4056 = 4'h7 == lineCounter ? frameBuffer_7_117 : _GEN_4055; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4057 = 4'h8 == lineCounter ? frameBuffer_8_117 : _GEN_4056; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4058 = 4'h9 == lineCounter ? frameBuffer_9_117 : _GEN_4057; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4059 = 4'ha == lineCounter ? frameBuffer_10_117 : _GEN_4058; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4060 = 4'hb == lineCounter ? frameBuffer_11_117 : _GEN_4059; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4061 = 4'hc == lineCounter ? frameBuffer_12_117 : _GEN_4060; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4062 = 4'hd == lineCounter ? frameBuffer_13_117 : _GEN_4061; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4063 = 4'he == lineCounter ? frameBuffer_14_117 : _GEN_4062; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4066 = 4'h1 == lineCounter ? frameBuffer_1_118 : frameBuffer_0_118; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4067 = 4'h2 == lineCounter ? frameBuffer_2_118 : _GEN_4066; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4068 = 4'h3 == lineCounter ? frameBuffer_3_118 : _GEN_4067; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4069 = 4'h4 == lineCounter ? frameBuffer_4_118 : _GEN_4068; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4070 = 4'h5 == lineCounter ? frameBuffer_5_118 : _GEN_4069; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4071 = 4'h6 == lineCounter ? frameBuffer_6_118 : _GEN_4070; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4072 = 4'h7 == lineCounter ? frameBuffer_7_118 : _GEN_4071; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4073 = 4'h8 == lineCounter ? frameBuffer_8_118 : _GEN_4072; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4074 = 4'h9 == lineCounter ? frameBuffer_9_118 : _GEN_4073; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4075 = 4'ha == lineCounter ? frameBuffer_10_118 : _GEN_4074; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4076 = 4'hb == lineCounter ? frameBuffer_11_118 : _GEN_4075; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4077 = 4'hc == lineCounter ? frameBuffer_12_118 : _GEN_4076; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4078 = 4'hd == lineCounter ? frameBuffer_13_118 : _GEN_4077; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4079 = 4'he == lineCounter ? frameBuffer_14_118 : _GEN_4078; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4082 = 4'h1 == lineCounter ? frameBuffer_1_119 : frameBuffer_0_119; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4083 = 4'h2 == lineCounter ? frameBuffer_2_119 : _GEN_4082; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4084 = 4'h3 == lineCounter ? frameBuffer_3_119 : _GEN_4083; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4085 = 4'h4 == lineCounter ? frameBuffer_4_119 : _GEN_4084; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4086 = 4'h5 == lineCounter ? frameBuffer_5_119 : _GEN_4085; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4087 = 4'h6 == lineCounter ? frameBuffer_6_119 : _GEN_4086; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4088 = 4'h7 == lineCounter ? frameBuffer_7_119 : _GEN_4087; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4089 = 4'h8 == lineCounter ? frameBuffer_8_119 : _GEN_4088; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4090 = 4'h9 == lineCounter ? frameBuffer_9_119 : _GEN_4089; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4091 = 4'ha == lineCounter ? frameBuffer_10_119 : _GEN_4090; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4092 = 4'hb == lineCounter ? frameBuffer_11_119 : _GEN_4091; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4093 = 4'hc == lineCounter ? frameBuffer_12_119 : _GEN_4092; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4094 = 4'hd == lineCounter ? frameBuffer_13_119 : _GEN_4093; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4095 = 4'he == lineCounter ? frameBuffer_14_119 : _GEN_4094; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4098 = 4'h1 == lineCounter ? frameBuffer_1_120 : frameBuffer_0_120; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4099 = 4'h2 == lineCounter ? frameBuffer_2_120 : _GEN_4098; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4100 = 4'h3 == lineCounter ? frameBuffer_3_120 : _GEN_4099; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4101 = 4'h4 == lineCounter ? frameBuffer_4_120 : _GEN_4100; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4102 = 4'h5 == lineCounter ? frameBuffer_5_120 : _GEN_4101; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4103 = 4'h6 == lineCounter ? frameBuffer_6_120 : _GEN_4102; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4104 = 4'h7 == lineCounter ? frameBuffer_7_120 : _GEN_4103; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4105 = 4'h8 == lineCounter ? frameBuffer_8_120 : _GEN_4104; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4106 = 4'h9 == lineCounter ? frameBuffer_9_120 : _GEN_4105; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4107 = 4'ha == lineCounter ? frameBuffer_10_120 : _GEN_4106; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4108 = 4'hb == lineCounter ? frameBuffer_11_120 : _GEN_4107; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4109 = 4'hc == lineCounter ? frameBuffer_12_120 : _GEN_4108; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4110 = 4'hd == lineCounter ? frameBuffer_13_120 : _GEN_4109; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4111 = 4'he == lineCounter ? frameBuffer_14_120 : _GEN_4110; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4114 = 4'h1 == lineCounter ? frameBuffer_1_121 : frameBuffer_0_121; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4115 = 4'h2 == lineCounter ? frameBuffer_2_121 : _GEN_4114; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4116 = 4'h3 == lineCounter ? frameBuffer_3_121 : _GEN_4115; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4117 = 4'h4 == lineCounter ? frameBuffer_4_121 : _GEN_4116; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4118 = 4'h5 == lineCounter ? frameBuffer_5_121 : _GEN_4117; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4119 = 4'h6 == lineCounter ? frameBuffer_6_121 : _GEN_4118; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4120 = 4'h7 == lineCounter ? frameBuffer_7_121 : _GEN_4119; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4121 = 4'h8 == lineCounter ? frameBuffer_8_121 : _GEN_4120; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4122 = 4'h9 == lineCounter ? frameBuffer_9_121 : _GEN_4121; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4123 = 4'ha == lineCounter ? frameBuffer_10_121 : _GEN_4122; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4124 = 4'hb == lineCounter ? frameBuffer_11_121 : _GEN_4123; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4125 = 4'hc == lineCounter ? frameBuffer_12_121 : _GEN_4124; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4126 = 4'hd == lineCounter ? frameBuffer_13_121 : _GEN_4125; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4127 = 4'he == lineCounter ? frameBuffer_14_121 : _GEN_4126; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4130 = 4'h1 == lineCounter ? frameBuffer_1_122 : frameBuffer_0_122; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4131 = 4'h2 == lineCounter ? frameBuffer_2_122 : _GEN_4130; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4132 = 4'h3 == lineCounter ? frameBuffer_3_122 : _GEN_4131; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4133 = 4'h4 == lineCounter ? frameBuffer_4_122 : _GEN_4132; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4134 = 4'h5 == lineCounter ? frameBuffer_5_122 : _GEN_4133; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4135 = 4'h6 == lineCounter ? frameBuffer_6_122 : _GEN_4134; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4136 = 4'h7 == lineCounter ? frameBuffer_7_122 : _GEN_4135; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4137 = 4'h8 == lineCounter ? frameBuffer_8_122 : _GEN_4136; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4138 = 4'h9 == lineCounter ? frameBuffer_9_122 : _GEN_4137; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4139 = 4'ha == lineCounter ? frameBuffer_10_122 : _GEN_4138; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4140 = 4'hb == lineCounter ? frameBuffer_11_122 : _GEN_4139; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4141 = 4'hc == lineCounter ? frameBuffer_12_122 : _GEN_4140; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4142 = 4'hd == lineCounter ? frameBuffer_13_122 : _GEN_4141; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4143 = 4'he == lineCounter ? frameBuffer_14_122 : _GEN_4142; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4146 = 4'h1 == lineCounter ? frameBuffer_1_123 : frameBuffer_0_123; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4147 = 4'h2 == lineCounter ? frameBuffer_2_123 : _GEN_4146; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4148 = 4'h3 == lineCounter ? frameBuffer_3_123 : _GEN_4147; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4149 = 4'h4 == lineCounter ? frameBuffer_4_123 : _GEN_4148; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4150 = 4'h5 == lineCounter ? frameBuffer_5_123 : _GEN_4149; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4151 = 4'h6 == lineCounter ? frameBuffer_6_123 : _GEN_4150; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4152 = 4'h7 == lineCounter ? frameBuffer_7_123 : _GEN_4151; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4153 = 4'h8 == lineCounter ? frameBuffer_8_123 : _GEN_4152; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4154 = 4'h9 == lineCounter ? frameBuffer_9_123 : _GEN_4153; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4155 = 4'ha == lineCounter ? frameBuffer_10_123 : _GEN_4154; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4156 = 4'hb == lineCounter ? frameBuffer_11_123 : _GEN_4155; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4157 = 4'hc == lineCounter ? frameBuffer_12_123 : _GEN_4156; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4158 = 4'hd == lineCounter ? frameBuffer_13_123 : _GEN_4157; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4159 = 4'he == lineCounter ? frameBuffer_14_123 : _GEN_4158; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4162 = 4'h1 == lineCounter ? frameBuffer_1_124 : frameBuffer_0_124; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4163 = 4'h2 == lineCounter ? frameBuffer_2_124 : _GEN_4162; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4164 = 4'h3 == lineCounter ? frameBuffer_3_124 : _GEN_4163; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4165 = 4'h4 == lineCounter ? frameBuffer_4_124 : _GEN_4164; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4166 = 4'h5 == lineCounter ? frameBuffer_5_124 : _GEN_4165; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4167 = 4'h6 == lineCounter ? frameBuffer_6_124 : _GEN_4166; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4168 = 4'h7 == lineCounter ? frameBuffer_7_124 : _GEN_4167; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4169 = 4'h8 == lineCounter ? frameBuffer_8_124 : _GEN_4168; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4170 = 4'h9 == lineCounter ? frameBuffer_9_124 : _GEN_4169; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4171 = 4'ha == lineCounter ? frameBuffer_10_124 : _GEN_4170; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4172 = 4'hb == lineCounter ? frameBuffer_11_124 : _GEN_4171; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4173 = 4'hc == lineCounter ? frameBuffer_12_124 : _GEN_4172; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4174 = 4'hd == lineCounter ? frameBuffer_13_124 : _GEN_4173; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4175 = 4'he == lineCounter ? frameBuffer_14_124 : _GEN_4174; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4178 = 4'h1 == lineCounter ? frameBuffer_1_125 : frameBuffer_0_125; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4179 = 4'h2 == lineCounter ? frameBuffer_2_125 : _GEN_4178; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4180 = 4'h3 == lineCounter ? frameBuffer_3_125 : _GEN_4179; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4181 = 4'h4 == lineCounter ? frameBuffer_4_125 : _GEN_4180; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4182 = 4'h5 == lineCounter ? frameBuffer_5_125 : _GEN_4181; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4183 = 4'h6 == lineCounter ? frameBuffer_6_125 : _GEN_4182; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4184 = 4'h7 == lineCounter ? frameBuffer_7_125 : _GEN_4183; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4185 = 4'h8 == lineCounter ? frameBuffer_8_125 : _GEN_4184; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4186 = 4'h9 == lineCounter ? frameBuffer_9_125 : _GEN_4185; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4187 = 4'ha == lineCounter ? frameBuffer_10_125 : _GEN_4186; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4188 = 4'hb == lineCounter ? frameBuffer_11_125 : _GEN_4187; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4189 = 4'hc == lineCounter ? frameBuffer_12_125 : _GEN_4188; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4190 = 4'hd == lineCounter ? frameBuffer_13_125 : _GEN_4189; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4191 = 4'he == lineCounter ? frameBuffer_14_125 : _GEN_4190; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4194 = 4'h1 == lineCounter ? frameBuffer_1_126 : frameBuffer_0_126; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4195 = 4'h2 == lineCounter ? frameBuffer_2_126 : _GEN_4194; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4196 = 4'h3 == lineCounter ? frameBuffer_3_126 : _GEN_4195; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4197 = 4'h4 == lineCounter ? frameBuffer_4_126 : _GEN_4196; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4198 = 4'h5 == lineCounter ? frameBuffer_5_126 : _GEN_4197; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4199 = 4'h6 == lineCounter ? frameBuffer_6_126 : _GEN_4198; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4200 = 4'h7 == lineCounter ? frameBuffer_7_126 : _GEN_4199; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4201 = 4'h8 == lineCounter ? frameBuffer_8_126 : _GEN_4200; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4202 = 4'h9 == lineCounter ? frameBuffer_9_126 : _GEN_4201; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4203 = 4'ha == lineCounter ? frameBuffer_10_126 : _GEN_4202; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4204 = 4'hb == lineCounter ? frameBuffer_11_126 : _GEN_4203; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4205 = 4'hc == lineCounter ? frameBuffer_12_126 : _GEN_4204; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4206 = 4'hd == lineCounter ? frameBuffer_13_126 : _GEN_4205; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4207 = 4'he == lineCounter ? frameBuffer_14_126 : _GEN_4206; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4210 = 4'h1 == lineCounter ? frameBuffer_1_127 : frameBuffer_0_127; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4211 = 4'h2 == lineCounter ? frameBuffer_2_127 : _GEN_4210; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4212 = 4'h3 == lineCounter ? frameBuffer_3_127 : _GEN_4211; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4213 = 4'h4 == lineCounter ? frameBuffer_4_127 : _GEN_4212; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4214 = 4'h5 == lineCounter ? frameBuffer_5_127 : _GEN_4213; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4215 = 4'h6 == lineCounter ? frameBuffer_6_127 : _GEN_4214; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4216 = 4'h7 == lineCounter ? frameBuffer_7_127 : _GEN_4215; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4217 = 4'h8 == lineCounter ? frameBuffer_8_127 : _GEN_4216; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4218 = 4'h9 == lineCounter ? frameBuffer_9_127 : _GEN_4217; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4219 = 4'ha == lineCounter ? frameBuffer_10_127 : _GEN_4218; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4220 = 4'hb == lineCounter ? frameBuffer_11_127 : _GEN_4219; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4221 = 4'hc == lineCounter ? frameBuffer_12_127 : _GEN_4220; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4222 = 4'hd == lineCounter ? frameBuffer_13_127 : _GEN_4221; // @[BufferAMSNew.scala 67:{15,15}]
  wire [7:0] _GEN_4223 = 4'he == lineCounter ? frameBuffer_14_127 : _GEN_4222; // @[BufferAMSNew.scala 67:{15,15}]
  wire [16:0] _GEN_4353 = reset ? 17'h0 : _GEN_2161; // @[BufferAMSNew.scala 14:{33,33}]
  wire [16:0] _GEN_4354 = reset ? 17'h0 : _GEN_2162; // @[BufferAMSNew.scala 14:{33,33}]
  wire [16:0] _GEN_4355 = reset ? 17'h0 : _GEN_2163; // @[BufferAMSNew.scala 14:{33,33}]
  wire [16:0] _GEN_4356 = reset ? 17'h0 : _GEN_2164; // @[BufferAMSNew.scala 14:{33,33}]
  wire [16:0] _GEN_4357 = reset ? 17'h0 : _GEN_2165; // @[BufferAMSNew.scala 14:{33,33}]
  wire [16:0] _GEN_4358 = reset ? 17'h0 : _GEN_2166; // @[BufferAMSNew.scala 14:{33,33}]
  wire [16:0] _GEN_4359 = reset ? 17'h0 : _GEN_2167; // @[BufferAMSNew.scala 14:{33,33}]
  wire [16:0] _GEN_4360 = reset ? 17'h0 : _GEN_2168; // @[BufferAMSNew.scala 14:{33,33}]
  assign io_zeroSums_0 = zeroAccumulators_0; // @[BufferAMSNew.scala 63:15]
  assign io_zeroSums_1 = zeroAccumulators_1; // @[BufferAMSNew.scala 63:15]
  assign io_zeroSums_2 = zeroAccumulators_2; // @[BufferAMSNew.scala 63:15]
  assign io_zeroSums_3 = zeroAccumulators_3; // @[BufferAMSNew.scala 63:15]
  assign io_zeroSums_4 = zeroAccumulators_4; // @[BufferAMSNew.scala 63:15]
  assign io_zeroSums_5 = zeroAccumulators_5; // @[BufferAMSNew.scala 63:15]
  assign io_zeroSums_6 = zeroAccumulators_6; // @[BufferAMSNew.scala 63:15]
  assign io_zeroSums_7 = zeroAccumulators_7; // @[BufferAMSNew.scala 63:15]
  assign io_indicesOut_0 = indexAccumulators_0; // @[BufferAMSNew.scala 64:17]
  assign io_indicesOut_1 = indexAccumulators_1; // @[BufferAMSNew.scala 64:17]
  assign io_indicesOut_2 = indexAccumulators_2; // @[BufferAMSNew.scala 64:17]
  assign io_indicesOut_3 = indexAccumulators_3; // @[BufferAMSNew.scala 64:17]
  assign io_indicesOut_4 = indexAccumulators_4; // @[BufferAMSNew.scala 64:17]
  assign io_indicesOut_5 = indexAccumulators_5; // @[BufferAMSNew.scala 64:17]
  assign io_indicesOut_6 = indexAccumulators_6; // @[BufferAMSNew.scala 64:17]
  assign io_indicesOut_7 = indexAccumulators_7; // @[BufferAMSNew.scala 64:17]
  assign io_frameOut_0 = 4'hf == lineCounter ? frameBuffer_15_0 : _GEN_2191; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_1 = 4'hf == lineCounter ? frameBuffer_15_1 : _GEN_2207; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_2 = 4'hf == lineCounter ? frameBuffer_15_2 : _GEN_2223; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_3 = 4'hf == lineCounter ? frameBuffer_15_3 : _GEN_2239; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_4 = 4'hf == lineCounter ? frameBuffer_15_4 : _GEN_2255; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_5 = 4'hf == lineCounter ? frameBuffer_15_5 : _GEN_2271; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_6 = 4'hf == lineCounter ? frameBuffer_15_6 : _GEN_2287; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_7 = 4'hf == lineCounter ? frameBuffer_15_7 : _GEN_2303; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_8 = 4'hf == lineCounter ? frameBuffer_15_8 : _GEN_2319; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_9 = 4'hf == lineCounter ? frameBuffer_15_9 : _GEN_2335; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_10 = 4'hf == lineCounter ? frameBuffer_15_10 : _GEN_2351; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_11 = 4'hf == lineCounter ? frameBuffer_15_11 : _GEN_2367; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_12 = 4'hf == lineCounter ? frameBuffer_15_12 : _GEN_2383; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_13 = 4'hf == lineCounter ? frameBuffer_15_13 : _GEN_2399; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_14 = 4'hf == lineCounter ? frameBuffer_15_14 : _GEN_2415; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_15 = 4'hf == lineCounter ? frameBuffer_15_15 : _GEN_2431; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_16 = 4'hf == lineCounter ? frameBuffer_15_16 : _GEN_2447; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_17 = 4'hf == lineCounter ? frameBuffer_15_17 : _GEN_2463; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_18 = 4'hf == lineCounter ? frameBuffer_15_18 : _GEN_2479; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_19 = 4'hf == lineCounter ? frameBuffer_15_19 : _GEN_2495; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_20 = 4'hf == lineCounter ? frameBuffer_15_20 : _GEN_2511; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_21 = 4'hf == lineCounter ? frameBuffer_15_21 : _GEN_2527; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_22 = 4'hf == lineCounter ? frameBuffer_15_22 : _GEN_2543; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_23 = 4'hf == lineCounter ? frameBuffer_15_23 : _GEN_2559; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_24 = 4'hf == lineCounter ? frameBuffer_15_24 : _GEN_2575; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_25 = 4'hf == lineCounter ? frameBuffer_15_25 : _GEN_2591; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_26 = 4'hf == lineCounter ? frameBuffer_15_26 : _GEN_2607; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_27 = 4'hf == lineCounter ? frameBuffer_15_27 : _GEN_2623; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_28 = 4'hf == lineCounter ? frameBuffer_15_28 : _GEN_2639; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_29 = 4'hf == lineCounter ? frameBuffer_15_29 : _GEN_2655; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_30 = 4'hf == lineCounter ? frameBuffer_15_30 : _GEN_2671; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_31 = 4'hf == lineCounter ? frameBuffer_15_31 : _GEN_2687; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_32 = 4'hf == lineCounter ? frameBuffer_15_32 : _GEN_2703; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_33 = 4'hf == lineCounter ? frameBuffer_15_33 : _GEN_2719; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_34 = 4'hf == lineCounter ? frameBuffer_15_34 : _GEN_2735; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_35 = 4'hf == lineCounter ? frameBuffer_15_35 : _GEN_2751; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_36 = 4'hf == lineCounter ? frameBuffer_15_36 : _GEN_2767; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_37 = 4'hf == lineCounter ? frameBuffer_15_37 : _GEN_2783; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_38 = 4'hf == lineCounter ? frameBuffer_15_38 : _GEN_2799; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_39 = 4'hf == lineCounter ? frameBuffer_15_39 : _GEN_2815; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_40 = 4'hf == lineCounter ? frameBuffer_15_40 : _GEN_2831; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_41 = 4'hf == lineCounter ? frameBuffer_15_41 : _GEN_2847; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_42 = 4'hf == lineCounter ? frameBuffer_15_42 : _GEN_2863; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_43 = 4'hf == lineCounter ? frameBuffer_15_43 : _GEN_2879; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_44 = 4'hf == lineCounter ? frameBuffer_15_44 : _GEN_2895; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_45 = 4'hf == lineCounter ? frameBuffer_15_45 : _GEN_2911; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_46 = 4'hf == lineCounter ? frameBuffer_15_46 : _GEN_2927; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_47 = 4'hf == lineCounter ? frameBuffer_15_47 : _GEN_2943; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_48 = 4'hf == lineCounter ? frameBuffer_15_48 : _GEN_2959; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_49 = 4'hf == lineCounter ? frameBuffer_15_49 : _GEN_2975; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_50 = 4'hf == lineCounter ? frameBuffer_15_50 : _GEN_2991; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_51 = 4'hf == lineCounter ? frameBuffer_15_51 : _GEN_3007; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_52 = 4'hf == lineCounter ? frameBuffer_15_52 : _GEN_3023; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_53 = 4'hf == lineCounter ? frameBuffer_15_53 : _GEN_3039; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_54 = 4'hf == lineCounter ? frameBuffer_15_54 : _GEN_3055; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_55 = 4'hf == lineCounter ? frameBuffer_15_55 : _GEN_3071; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_56 = 4'hf == lineCounter ? frameBuffer_15_56 : _GEN_3087; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_57 = 4'hf == lineCounter ? frameBuffer_15_57 : _GEN_3103; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_58 = 4'hf == lineCounter ? frameBuffer_15_58 : _GEN_3119; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_59 = 4'hf == lineCounter ? frameBuffer_15_59 : _GEN_3135; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_60 = 4'hf == lineCounter ? frameBuffer_15_60 : _GEN_3151; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_61 = 4'hf == lineCounter ? frameBuffer_15_61 : _GEN_3167; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_62 = 4'hf == lineCounter ? frameBuffer_15_62 : _GEN_3183; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_63 = 4'hf == lineCounter ? frameBuffer_15_63 : _GEN_3199; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_64 = 4'hf == lineCounter ? frameBuffer_15_64 : _GEN_3215; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_65 = 4'hf == lineCounter ? frameBuffer_15_65 : _GEN_3231; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_66 = 4'hf == lineCounter ? frameBuffer_15_66 : _GEN_3247; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_67 = 4'hf == lineCounter ? frameBuffer_15_67 : _GEN_3263; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_68 = 4'hf == lineCounter ? frameBuffer_15_68 : _GEN_3279; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_69 = 4'hf == lineCounter ? frameBuffer_15_69 : _GEN_3295; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_70 = 4'hf == lineCounter ? frameBuffer_15_70 : _GEN_3311; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_71 = 4'hf == lineCounter ? frameBuffer_15_71 : _GEN_3327; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_72 = 4'hf == lineCounter ? frameBuffer_15_72 : _GEN_3343; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_73 = 4'hf == lineCounter ? frameBuffer_15_73 : _GEN_3359; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_74 = 4'hf == lineCounter ? frameBuffer_15_74 : _GEN_3375; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_75 = 4'hf == lineCounter ? frameBuffer_15_75 : _GEN_3391; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_76 = 4'hf == lineCounter ? frameBuffer_15_76 : _GEN_3407; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_77 = 4'hf == lineCounter ? frameBuffer_15_77 : _GEN_3423; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_78 = 4'hf == lineCounter ? frameBuffer_15_78 : _GEN_3439; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_79 = 4'hf == lineCounter ? frameBuffer_15_79 : _GEN_3455; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_80 = 4'hf == lineCounter ? frameBuffer_15_80 : _GEN_3471; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_81 = 4'hf == lineCounter ? frameBuffer_15_81 : _GEN_3487; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_82 = 4'hf == lineCounter ? frameBuffer_15_82 : _GEN_3503; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_83 = 4'hf == lineCounter ? frameBuffer_15_83 : _GEN_3519; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_84 = 4'hf == lineCounter ? frameBuffer_15_84 : _GEN_3535; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_85 = 4'hf == lineCounter ? frameBuffer_15_85 : _GEN_3551; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_86 = 4'hf == lineCounter ? frameBuffer_15_86 : _GEN_3567; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_87 = 4'hf == lineCounter ? frameBuffer_15_87 : _GEN_3583; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_88 = 4'hf == lineCounter ? frameBuffer_15_88 : _GEN_3599; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_89 = 4'hf == lineCounter ? frameBuffer_15_89 : _GEN_3615; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_90 = 4'hf == lineCounter ? frameBuffer_15_90 : _GEN_3631; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_91 = 4'hf == lineCounter ? frameBuffer_15_91 : _GEN_3647; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_92 = 4'hf == lineCounter ? frameBuffer_15_92 : _GEN_3663; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_93 = 4'hf == lineCounter ? frameBuffer_15_93 : _GEN_3679; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_94 = 4'hf == lineCounter ? frameBuffer_15_94 : _GEN_3695; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_95 = 4'hf == lineCounter ? frameBuffer_15_95 : _GEN_3711; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_96 = 4'hf == lineCounter ? frameBuffer_15_96 : _GEN_3727; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_97 = 4'hf == lineCounter ? frameBuffer_15_97 : _GEN_3743; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_98 = 4'hf == lineCounter ? frameBuffer_15_98 : _GEN_3759; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_99 = 4'hf == lineCounter ? frameBuffer_15_99 : _GEN_3775; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_100 = 4'hf == lineCounter ? frameBuffer_15_100 : _GEN_3791; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_101 = 4'hf == lineCounter ? frameBuffer_15_101 : _GEN_3807; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_102 = 4'hf == lineCounter ? frameBuffer_15_102 : _GEN_3823; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_103 = 4'hf == lineCounter ? frameBuffer_15_103 : _GEN_3839; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_104 = 4'hf == lineCounter ? frameBuffer_15_104 : _GEN_3855; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_105 = 4'hf == lineCounter ? frameBuffer_15_105 : _GEN_3871; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_106 = 4'hf == lineCounter ? frameBuffer_15_106 : _GEN_3887; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_107 = 4'hf == lineCounter ? frameBuffer_15_107 : _GEN_3903; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_108 = 4'hf == lineCounter ? frameBuffer_15_108 : _GEN_3919; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_109 = 4'hf == lineCounter ? frameBuffer_15_109 : _GEN_3935; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_110 = 4'hf == lineCounter ? frameBuffer_15_110 : _GEN_3951; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_111 = 4'hf == lineCounter ? frameBuffer_15_111 : _GEN_3967; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_112 = 4'hf == lineCounter ? frameBuffer_15_112 : _GEN_3983; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_113 = 4'hf == lineCounter ? frameBuffer_15_113 : _GEN_3999; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_114 = 4'hf == lineCounter ? frameBuffer_15_114 : _GEN_4015; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_115 = 4'hf == lineCounter ? frameBuffer_15_115 : _GEN_4031; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_116 = 4'hf == lineCounter ? frameBuffer_15_116 : _GEN_4047; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_117 = 4'hf == lineCounter ? frameBuffer_15_117 : _GEN_4063; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_118 = 4'hf == lineCounter ? frameBuffer_15_118 : _GEN_4079; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_119 = 4'hf == lineCounter ? frameBuffer_15_119 : _GEN_4095; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_120 = 4'hf == lineCounter ? frameBuffer_15_120 : _GEN_4111; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_121 = 4'hf == lineCounter ? frameBuffer_15_121 : _GEN_4127; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_122 = 4'hf == lineCounter ? frameBuffer_15_122 : _GEN_4143; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_123 = 4'hf == lineCounter ? frameBuffer_15_123 : _GEN_4159; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_124 = 4'hf == lineCounter ? frameBuffer_15_124 : _GEN_4175; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_125 = 4'hf == lineCounter ? frameBuffer_15_125 : _GEN_4191; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_126 = 4'hf == lineCounter ? frameBuffer_15_126 : _GEN_4207; // @[BufferAMSNew.scala 67:{15,15}]
  assign io_frameOut_127 = 4'hf == lineCounter ? frameBuffer_15_127 : _GEN_4223; // @[BufferAMSNew.scala 67:{15,15}]
  always @(posedge clock) begin
    zeroAccumulators_0 <= _GEN_4353[7:0]; // @[BufferAMSNew.scala 14:{33,33}]
    zeroAccumulators_1 <= _GEN_4354[7:0]; // @[BufferAMSNew.scala 14:{33,33}]
    zeroAccumulators_2 <= _GEN_4355[7:0]; // @[BufferAMSNew.scala 14:{33,33}]
    zeroAccumulators_3 <= _GEN_4356[7:0]; // @[BufferAMSNew.scala 14:{33,33}]
    zeroAccumulators_4 <= _GEN_4357[7:0]; // @[BufferAMSNew.scala 14:{33,33}]
    zeroAccumulators_5 <= _GEN_4358[7:0]; // @[BufferAMSNew.scala 14:{33,33}]
    zeroAccumulators_6 <= _GEN_4359[7:0]; // @[BufferAMSNew.scala 14:{33,33}]
    zeroAccumulators_7 <= _GEN_4360[7:0]; // @[BufferAMSNew.scala 14:{33,33}]
    if (reset) begin // @[BufferAMSNew.scala 17:34]
      indexAccumulators_0 <= 4'h0; // @[BufferAMSNew.scala 17:34]
    end else if (lineCounter == 4'hf) begin // @[BufferAMSNew.scala 28:30]
      indexAccumulators_0 <= 4'h0; // @[BufferAMSNew.scala 31:23]
    end else if (zeroAccumulators_0 < zeroAccumulators_1) begin // @[BufferAMSNew.scala 47:61]
      indexAccumulators_0 <= indexAccumulators_1; // @[BufferAMSNew.scala 55:32]
    end else if (zeroAccumulators_0 < zeroAccumulators_1) begin // @[BufferAMSNew.scala 47:61]
      indexAccumulators_0 <= indexAccumulators_1; // @[BufferAMSNew.scala 55:32]
    end else begin
      indexAccumulators_0 <= _GEN_2138;
    end
    if (reset) begin // @[BufferAMSNew.scala 17:34]
      indexAccumulators_1 <= 4'h1; // @[BufferAMSNew.scala 17:34]
    end else if (lineCounter == 4'hf) begin // @[BufferAMSNew.scala 28:30]
      indexAccumulators_1 <= 4'h1; // @[BufferAMSNew.scala 31:23]
    end else if (zeroAccumulators_0 < zeroAccumulators_1) begin // @[BufferAMSNew.scala 47:61]
      indexAccumulators_1 <= indexAccumulators_0; // @[BufferAMSNew.scala 56:36]
    end else if (zeroAccumulators_1 < zeroAccumulators_2) begin // @[BufferAMSNew.scala 47:61]
      indexAccumulators_1 <= indexAccumulators_2; // @[BufferAMSNew.scala 55:32]
    end else begin
      indexAccumulators_1 <= _GEN_2151;
    end
    if (reset) begin // @[BufferAMSNew.scala 17:34]
      indexAccumulators_2 <= 4'h2; // @[BufferAMSNew.scala 17:34]
    end else if (lineCounter == 4'hf) begin // @[BufferAMSNew.scala 28:30]
      indexAccumulators_2 <= 4'h2; // @[BufferAMSNew.scala 31:23]
    end else if (zeroAccumulators_1 < zeroAccumulators_2) begin // @[BufferAMSNew.scala 47:61]
      indexAccumulators_2 <= indexAccumulators_1; // @[BufferAMSNew.scala 56:36]
    end else if (zeroAccumulators_2 < zeroAccumulators_3) begin // @[BufferAMSNew.scala 47:61]
      indexAccumulators_2 <= indexAccumulators_3; // @[BufferAMSNew.scala 55:32]
    end else begin
      indexAccumulators_2 <= _GEN_2143;
    end
    if (reset) begin // @[BufferAMSNew.scala 17:34]
      indexAccumulators_3 <= 4'h3; // @[BufferAMSNew.scala 17:34]
    end else if (lineCounter == 4'hf) begin // @[BufferAMSNew.scala 28:30]
      indexAccumulators_3 <= 4'h3; // @[BufferAMSNew.scala 31:23]
    end else if (zeroAccumulators_2 < zeroAccumulators_3) begin // @[BufferAMSNew.scala 47:61]
      indexAccumulators_3 <= indexAccumulators_2; // @[BufferAMSNew.scala 56:36]
    end else if (zeroAccumulators_3 < zeroAccumulators_4) begin // @[BufferAMSNew.scala 47:61]
      indexAccumulators_3 <= indexAccumulators_4; // @[BufferAMSNew.scala 55:32]
    end else begin
      indexAccumulators_3 <= _GEN_2131;
    end
    if (reset) begin // @[BufferAMSNew.scala 17:34]
      indexAccumulators_4 <= 4'h4; // @[BufferAMSNew.scala 17:34]
    end else if (lineCounter == 4'hf) begin // @[BufferAMSNew.scala 28:30]
      indexAccumulators_4 <= 4'h4; // @[BufferAMSNew.scala 31:23]
    end else if (zeroAccumulators_3 < zeroAccumulators_4) begin // @[BufferAMSNew.scala 47:61]
      indexAccumulators_4 <= indexAccumulators_3; // @[BufferAMSNew.scala 56:36]
    end else if (zeroAccumulators_4 < zeroAccumulators_5) begin // @[BufferAMSNew.scala 47:61]
      indexAccumulators_4 <= indexAccumulators_5; // @[BufferAMSNew.scala 55:32]
    end else begin
      indexAccumulators_4 <= _GEN_2115;
    end
    if (reset) begin // @[BufferAMSNew.scala 17:34]
      indexAccumulators_5 <= 4'h5; // @[BufferAMSNew.scala 17:34]
    end else if (lineCounter == 4'hf) begin // @[BufferAMSNew.scala 28:30]
      indexAccumulators_5 <= 4'h5; // @[BufferAMSNew.scala 31:23]
    end else if (zeroAccumulators_4 < zeroAccumulators_5) begin // @[BufferAMSNew.scala 47:61]
      indexAccumulators_5 <= indexAccumulators_4; // @[BufferAMSNew.scala 56:36]
    end else if (zeroAccumulators_5 < zeroAccumulators_6) begin // @[BufferAMSNew.scala 47:61]
      indexAccumulators_5 <= indexAccumulators_6; // @[BufferAMSNew.scala 55:32]
    end else begin
      indexAccumulators_5 <= _GEN_2095;
    end
    if (reset) begin // @[BufferAMSNew.scala 17:34]
      indexAccumulators_6 <= 4'h6; // @[BufferAMSNew.scala 17:34]
    end else if (lineCounter == 4'hf) begin // @[BufferAMSNew.scala 28:30]
      indexAccumulators_6 <= 4'h6; // @[BufferAMSNew.scala 31:23]
    end else if (zeroAccumulators_5 < zeroAccumulators_6) begin // @[BufferAMSNew.scala 47:61]
      indexAccumulators_6 <= indexAccumulators_5; // @[BufferAMSNew.scala 56:36]
    end else if (zeroAccumulators_6 < zeroAccumulators_7) begin // @[BufferAMSNew.scala 47:61]
      indexAccumulators_6 <= indexAccumulators_7; // @[BufferAMSNew.scala 55:32]
    end else begin
      indexAccumulators_6 <= _GEN_2071;
    end
    if (reset) begin // @[BufferAMSNew.scala 17:34]
      indexAccumulators_7 <= 4'h7; // @[BufferAMSNew.scala 17:34]
    end else if (lineCounter == 4'hf) begin // @[BufferAMSNew.scala 28:30]
      indexAccumulators_7 <= 4'h7; // @[BufferAMSNew.scala 31:23]
    end else if (zeroAccumulators_6 < zeroAccumulators_7) begin // @[BufferAMSNew.scala 47:61]
      indexAccumulators_7 <= indexAccumulators_6; // @[BufferAMSNew.scala 56:36]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_0 <= io_adcValues_0; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_1 <= io_adcValues_1; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_2 <= io_adcValues_2; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_3 <= io_adcValues_3; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_4 <= io_adcValues_4; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_5 <= io_adcValues_5; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_6 <= io_adcValues_6; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_7 <= io_adcValues_7; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_8 <= io_adcValues_8; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_9 <= io_adcValues_9; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_10 <= io_adcValues_10; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_11 <= io_adcValues_11; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_12 <= io_adcValues_12; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_13 <= io_adcValues_13; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_14 <= io_adcValues_14; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_15 <= io_adcValues_15; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_16 <= io_adcValues_16; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_17 <= io_adcValues_17; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_18 <= io_adcValues_18; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_19 <= io_adcValues_19; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_20 <= io_adcValues_20; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_21 <= io_adcValues_21; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_22 <= io_adcValues_22; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_23 <= io_adcValues_23; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_24 <= io_adcValues_24; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_25 <= io_adcValues_25; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_26 <= io_adcValues_26; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_27 <= io_adcValues_27; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_28 <= io_adcValues_28; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_29 <= io_adcValues_29; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_30 <= io_adcValues_30; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_31 <= io_adcValues_31; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_32 <= io_adcValues_32; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_33 <= io_adcValues_33; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_34 <= io_adcValues_34; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_35 <= io_adcValues_35; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_36 <= io_adcValues_36; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_37 <= io_adcValues_37; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_38 <= io_adcValues_38; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_39 <= io_adcValues_39; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_40 <= io_adcValues_40; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_41 <= io_adcValues_41; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_42 <= io_adcValues_42; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_43 <= io_adcValues_43; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_44 <= io_adcValues_44; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_45 <= io_adcValues_45; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_46 <= io_adcValues_46; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_47 <= io_adcValues_47; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_48 <= io_adcValues_48; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_49 <= io_adcValues_49; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_50 <= io_adcValues_50; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_51 <= io_adcValues_51; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_52 <= io_adcValues_52; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_53 <= io_adcValues_53; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_54 <= io_adcValues_54; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_55 <= io_adcValues_55; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_56 <= io_adcValues_56; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_57 <= io_adcValues_57; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_58 <= io_adcValues_58; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_59 <= io_adcValues_59; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_60 <= io_adcValues_60; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_61 <= io_adcValues_61; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_62 <= io_adcValues_62; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_63 <= io_adcValues_63; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_64 <= io_adcValues_64; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_65 <= io_adcValues_65; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_66 <= io_adcValues_66; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_67 <= io_adcValues_67; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_68 <= io_adcValues_68; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_69 <= io_adcValues_69; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_70 <= io_adcValues_70; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_71 <= io_adcValues_71; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_72 <= io_adcValues_72; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_73 <= io_adcValues_73; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_74 <= io_adcValues_74; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_75 <= io_adcValues_75; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_76 <= io_adcValues_76; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_77 <= io_adcValues_77; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_78 <= io_adcValues_78; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_79 <= io_adcValues_79; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_80 <= io_adcValues_80; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_81 <= io_adcValues_81; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_82 <= io_adcValues_82; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_83 <= io_adcValues_83; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_84 <= io_adcValues_84; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_85 <= io_adcValues_85; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_86 <= io_adcValues_86; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_87 <= io_adcValues_87; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_88 <= io_adcValues_88; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_89 <= io_adcValues_89; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_90 <= io_adcValues_90; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_91 <= io_adcValues_91; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_92 <= io_adcValues_92; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_93 <= io_adcValues_93; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_94 <= io_adcValues_94; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_95 <= io_adcValues_95; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_96 <= io_adcValues_96; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_97 <= io_adcValues_97; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_98 <= io_adcValues_98; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_99 <= io_adcValues_99; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_100 <= io_adcValues_100; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_101 <= io_adcValues_101; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_102 <= io_adcValues_102; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_103 <= io_adcValues_103; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_104 <= io_adcValues_104; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_105 <= io_adcValues_105; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_106 <= io_adcValues_106; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_107 <= io_adcValues_107; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_108 <= io_adcValues_108; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_109 <= io_adcValues_109; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_110 <= io_adcValues_110; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_111 <= io_adcValues_111; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_112 <= io_adcValues_112; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_113 <= io_adcValues_113; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_114 <= io_adcValues_114; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_115 <= io_adcValues_115; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_116 <= io_adcValues_116; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_117 <= io_adcValues_117; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_118 <= io_adcValues_118; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_119 <= io_adcValues_119; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_120 <= io_adcValues_120; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_121 <= io_adcValues_121; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_122 <= io_adcValues_122; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_123 <= io_adcValues_123; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_124 <= io_adcValues_124; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_125 <= io_adcValues_125; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_126 <= io_adcValues_126; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h0 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_0_127 <= io_adcValues_127; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_0 <= io_adcValues_0; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_1 <= io_adcValues_1; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_2 <= io_adcValues_2; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_3 <= io_adcValues_3; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_4 <= io_adcValues_4; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_5 <= io_adcValues_5; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_6 <= io_adcValues_6; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_7 <= io_adcValues_7; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_8 <= io_adcValues_8; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_9 <= io_adcValues_9; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_10 <= io_adcValues_10; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_11 <= io_adcValues_11; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_12 <= io_adcValues_12; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_13 <= io_adcValues_13; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_14 <= io_adcValues_14; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_15 <= io_adcValues_15; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_16 <= io_adcValues_16; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_17 <= io_adcValues_17; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_18 <= io_adcValues_18; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_19 <= io_adcValues_19; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_20 <= io_adcValues_20; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_21 <= io_adcValues_21; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_22 <= io_adcValues_22; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_23 <= io_adcValues_23; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_24 <= io_adcValues_24; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_25 <= io_adcValues_25; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_26 <= io_adcValues_26; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_27 <= io_adcValues_27; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_28 <= io_adcValues_28; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_29 <= io_adcValues_29; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_30 <= io_adcValues_30; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_31 <= io_adcValues_31; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_32 <= io_adcValues_32; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_33 <= io_adcValues_33; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_34 <= io_adcValues_34; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_35 <= io_adcValues_35; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_36 <= io_adcValues_36; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_37 <= io_adcValues_37; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_38 <= io_adcValues_38; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_39 <= io_adcValues_39; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_40 <= io_adcValues_40; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_41 <= io_adcValues_41; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_42 <= io_adcValues_42; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_43 <= io_adcValues_43; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_44 <= io_adcValues_44; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_45 <= io_adcValues_45; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_46 <= io_adcValues_46; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_47 <= io_adcValues_47; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_48 <= io_adcValues_48; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_49 <= io_adcValues_49; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_50 <= io_adcValues_50; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_51 <= io_adcValues_51; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_52 <= io_adcValues_52; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_53 <= io_adcValues_53; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_54 <= io_adcValues_54; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_55 <= io_adcValues_55; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_56 <= io_adcValues_56; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_57 <= io_adcValues_57; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_58 <= io_adcValues_58; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_59 <= io_adcValues_59; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_60 <= io_adcValues_60; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_61 <= io_adcValues_61; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_62 <= io_adcValues_62; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_63 <= io_adcValues_63; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_64 <= io_adcValues_64; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_65 <= io_adcValues_65; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_66 <= io_adcValues_66; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_67 <= io_adcValues_67; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_68 <= io_adcValues_68; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_69 <= io_adcValues_69; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_70 <= io_adcValues_70; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_71 <= io_adcValues_71; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_72 <= io_adcValues_72; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_73 <= io_adcValues_73; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_74 <= io_adcValues_74; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_75 <= io_adcValues_75; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_76 <= io_adcValues_76; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_77 <= io_adcValues_77; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_78 <= io_adcValues_78; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_79 <= io_adcValues_79; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_80 <= io_adcValues_80; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_81 <= io_adcValues_81; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_82 <= io_adcValues_82; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_83 <= io_adcValues_83; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_84 <= io_adcValues_84; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_85 <= io_adcValues_85; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_86 <= io_adcValues_86; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_87 <= io_adcValues_87; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_88 <= io_adcValues_88; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_89 <= io_adcValues_89; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_90 <= io_adcValues_90; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_91 <= io_adcValues_91; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_92 <= io_adcValues_92; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_93 <= io_adcValues_93; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_94 <= io_adcValues_94; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_95 <= io_adcValues_95; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_96 <= io_adcValues_96; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_97 <= io_adcValues_97; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_98 <= io_adcValues_98; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_99 <= io_adcValues_99; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_100 <= io_adcValues_100; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_101 <= io_adcValues_101; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_102 <= io_adcValues_102; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_103 <= io_adcValues_103; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_104 <= io_adcValues_104; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_105 <= io_adcValues_105; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_106 <= io_adcValues_106; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_107 <= io_adcValues_107; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_108 <= io_adcValues_108; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_109 <= io_adcValues_109; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_110 <= io_adcValues_110; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_111 <= io_adcValues_111; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_112 <= io_adcValues_112; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_113 <= io_adcValues_113; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_114 <= io_adcValues_114; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_115 <= io_adcValues_115; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_116 <= io_adcValues_116; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_117 <= io_adcValues_117; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_118 <= io_adcValues_118; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_119 <= io_adcValues_119; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_120 <= io_adcValues_120; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_121 <= io_adcValues_121; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_122 <= io_adcValues_122; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_123 <= io_adcValues_123; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_124 <= io_adcValues_124; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_125 <= io_adcValues_125; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_126 <= io_adcValues_126; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h1 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_1_127 <= io_adcValues_127; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_0 <= io_adcValues_0; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_1 <= io_adcValues_1; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_2 <= io_adcValues_2; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_3 <= io_adcValues_3; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_4 <= io_adcValues_4; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_5 <= io_adcValues_5; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_6 <= io_adcValues_6; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_7 <= io_adcValues_7; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_8 <= io_adcValues_8; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_9 <= io_adcValues_9; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_10 <= io_adcValues_10; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_11 <= io_adcValues_11; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_12 <= io_adcValues_12; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_13 <= io_adcValues_13; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_14 <= io_adcValues_14; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_15 <= io_adcValues_15; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_16 <= io_adcValues_16; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_17 <= io_adcValues_17; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_18 <= io_adcValues_18; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_19 <= io_adcValues_19; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_20 <= io_adcValues_20; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_21 <= io_adcValues_21; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_22 <= io_adcValues_22; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_23 <= io_adcValues_23; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_24 <= io_adcValues_24; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_25 <= io_adcValues_25; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_26 <= io_adcValues_26; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_27 <= io_adcValues_27; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_28 <= io_adcValues_28; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_29 <= io_adcValues_29; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_30 <= io_adcValues_30; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_31 <= io_adcValues_31; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_32 <= io_adcValues_32; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_33 <= io_adcValues_33; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_34 <= io_adcValues_34; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_35 <= io_adcValues_35; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_36 <= io_adcValues_36; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_37 <= io_adcValues_37; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_38 <= io_adcValues_38; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_39 <= io_adcValues_39; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_40 <= io_adcValues_40; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_41 <= io_adcValues_41; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_42 <= io_adcValues_42; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_43 <= io_adcValues_43; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_44 <= io_adcValues_44; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_45 <= io_adcValues_45; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_46 <= io_adcValues_46; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_47 <= io_adcValues_47; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_48 <= io_adcValues_48; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_49 <= io_adcValues_49; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_50 <= io_adcValues_50; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_51 <= io_adcValues_51; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_52 <= io_adcValues_52; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_53 <= io_adcValues_53; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_54 <= io_adcValues_54; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_55 <= io_adcValues_55; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_56 <= io_adcValues_56; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_57 <= io_adcValues_57; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_58 <= io_adcValues_58; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_59 <= io_adcValues_59; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_60 <= io_adcValues_60; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_61 <= io_adcValues_61; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_62 <= io_adcValues_62; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_63 <= io_adcValues_63; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_64 <= io_adcValues_64; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_65 <= io_adcValues_65; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_66 <= io_adcValues_66; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_67 <= io_adcValues_67; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_68 <= io_adcValues_68; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_69 <= io_adcValues_69; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_70 <= io_adcValues_70; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_71 <= io_adcValues_71; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_72 <= io_adcValues_72; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_73 <= io_adcValues_73; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_74 <= io_adcValues_74; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_75 <= io_adcValues_75; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_76 <= io_adcValues_76; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_77 <= io_adcValues_77; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_78 <= io_adcValues_78; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_79 <= io_adcValues_79; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_80 <= io_adcValues_80; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_81 <= io_adcValues_81; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_82 <= io_adcValues_82; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_83 <= io_adcValues_83; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_84 <= io_adcValues_84; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_85 <= io_adcValues_85; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_86 <= io_adcValues_86; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_87 <= io_adcValues_87; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_88 <= io_adcValues_88; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_89 <= io_adcValues_89; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_90 <= io_adcValues_90; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_91 <= io_adcValues_91; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_92 <= io_adcValues_92; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_93 <= io_adcValues_93; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_94 <= io_adcValues_94; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_95 <= io_adcValues_95; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_96 <= io_adcValues_96; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_97 <= io_adcValues_97; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_98 <= io_adcValues_98; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_99 <= io_adcValues_99; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_100 <= io_adcValues_100; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_101 <= io_adcValues_101; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_102 <= io_adcValues_102; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_103 <= io_adcValues_103; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_104 <= io_adcValues_104; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_105 <= io_adcValues_105; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_106 <= io_adcValues_106; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_107 <= io_adcValues_107; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_108 <= io_adcValues_108; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_109 <= io_adcValues_109; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_110 <= io_adcValues_110; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_111 <= io_adcValues_111; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_112 <= io_adcValues_112; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_113 <= io_adcValues_113; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_114 <= io_adcValues_114; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_115 <= io_adcValues_115; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_116 <= io_adcValues_116; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_117 <= io_adcValues_117; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_118 <= io_adcValues_118; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_119 <= io_adcValues_119; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_120 <= io_adcValues_120; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_121 <= io_adcValues_121; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_122 <= io_adcValues_122; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_123 <= io_adcValues_123; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_124 <= io_adcValues_124; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_125 <= io_adcValues_125; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_126 <= io_adcValues_126; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h2 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_2_127 <= io_adcValues_127; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_0 <= io_adcValues_0; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_1 <= io_adcValues_1; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_2 <= io_adcValues_2; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_3 <= io_adcValues_3; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_4 <= io_adcValues_4; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_5 <= io_adcValues_5; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_6 <= io_adcValues_6; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_7 <= io_adcValues_7; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_8 <= io_adcValues_8; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_9 <= io_adcValues_9; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_10 <= io_adcValues_10; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_11 <= io_adcValues_11; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_12 <= io_adcValues_12; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_13 <= io_adcValues_13; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_14 <= io_adcValues_14; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_15 <= io_adcValues_15; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_16 <= io_adcValues_16; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_17 <= io_adcValues_17; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_18 <= io_adcValues_18; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_19 <= io_adcValues_19; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_20 <= io_adcValues_20; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_21 <= io_adcValues_21; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_22 <= io_adcValues_22; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_23 <= io_adcValues_23; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_24 <= io_adcValues_24; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_25 <= io_adcValues_25; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_26 <= io_adcValues_26; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_27 <= io_adcValues_27; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_28 <= io_adcValues_28; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_29 <= io_adcValues_29; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_30 <= io_adcValues_30; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_31 <= io_adcValues_31; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_32 <= io_adcValues_32; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_33 <= io_adcValues_33; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_34 <= io_adcValues_34; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_35 <= io_adcValues_35; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_36 <= io_adcValues_36; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_37 <= io_adcValues_37; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_38 <= io_adcValues_38; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_39 <= io_adcValues_39; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_40 <= io_adcValues_40; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_41 <= io_adcValues_41; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_42 <= io_adcValues_42; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_43 <= io_adcValues_43; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_44 <= io_adcValues_44; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_45 <= io_adcValues_45; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_46 <= io_adcValues_46; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_47 <= io_adcValues_47; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_48 <= io_adcValues_48; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_49 <= io_adcValues_49; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_50 <= io_adcValues_50; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_51 <= io_adcValues_51; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_52 <= io_adcValues_52; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_53 <= io_adcValues_53; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_54 <= io_adcValues_54; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_55 <= io_adcValues_55; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_56 <= io_adcValues_56; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_57 <= io_adcValues_57; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_58 <= io_adcValues_58; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_59 <= io_adcValues_59; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_60 <= io_adcValues_60; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_61 <= io_adcValues_61; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_62 <= io_adcValues_62; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_63 <= io_adcValues_63; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_64 <= io_adcValues_64; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_65 <= io_adcValues_65; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_66 <= io_adcValues_66; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_67 <= io_adcValues_67; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_68 <= io_adcValues_68; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_69 <= io_adcValues_69; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_70 <= io_adcValues_70; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_71 <= io_adcValues_71; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_72 <= io_adcValues_72; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_73 <= io_adcValues_73; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_74 <= io_adcValues_74; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_75 <= io_adcValues_75; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_76 <= io_adcValues_76; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_77 <= io_adcValues_77; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_78 <= io_adcValues_78; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_79 <= io_adcValues_79; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_80 <= io_adcValues_80; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_81 <= io_adcValues_81; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_82 <= io_adcValues_82; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_83 <= io_adcValues_83; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_84 <= io_adcValues_84; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_85 <= io_adcValues_85; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_86 <= io_adcValues_86; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_87 <= io_adcValues_87; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_88 <= io_adcValues_88; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_89 <= io_adcValues_89; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_90 <= io_adcValues_90; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_91 <= io_adcValues_91; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_92 <= io_adcValues_92; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_93 <= io_adcValues_93; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_94 <= io_adcValues_94; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_95 <= io_adcValues_95; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_96 <= io_adcValues_96; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_97 <= io_adcValues_97; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_98 <= io_adcValues_98; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_99 <= io_adcValues_99; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_100 <= io_adcValues_100; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_101 <= io_adcValues_101; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_102 <= io_adcValues_102; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_103 <= io_adcValues_103; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_104 <= io_adcValues_104; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_105 <= io_adcValues_105; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_106 <= io_adcValues_106; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_107 <= io_adcValues_107; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_108 <= io_adcValues_108; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_109 <= io_adcValues_109; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_110 <= io_adcValues_110; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_111 <= io_adcValues_111; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_112 <= io_adcValues_112; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_113 <= io_adcValues_113; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_114 <= io_adcValues_114; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_115 <= io_adcValues_115; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_116 <= io_adcValues_116; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_117 <= io_adcValues_117; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_118 <= io_adcValues_118; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_119 <= io_adcValues_119; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_120 <= io_adcValues_120; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_121 <= io_adcValues_121; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_122 <= io_adcValues_122; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_123 <= io_adcValues_123; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_124 <= io_adcValues_124; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_125 <= io_adcValues_125; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_126 <= io_adcValues_126; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h3 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_3_127 <= io_adcValues_127; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_0 <= io_adcValues_0; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_1 <= io_adcValues_1; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_2 <= io_adcValues_2; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_3 <= io_adcValues_3; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_4 <= io_adcValues_4; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_5 <= io_adcValues_5; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_6 <= io_adcValues_6; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_7 <= io_adcValues_7; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_8 <= io_adcValues_8; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_9 <= io_adcValues_9; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_10 <= io_adcValues_10; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_11 <= io_adcValues_11; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_12 <= io_adcValues_12; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_13 <= io_adcValues_13; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_14 <= io_adcValues_14; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_15 <= io_adcValues_15; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_16 <= io_adcValues_16; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_17 <= io_adcValues_17; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_18 <= io_adcValues_18; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_19 <= io_adcValues_19; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_20 <= io_adcValues_20; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_21 <= io_adcValues_21; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_22 <= io_adcValues_22; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_23 <= io_adcValues_23; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_24 <= io_adcValues_24; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_25 <= io_adcValues_25; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_26 <= io_adcValues_26; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_27 <= io_adcValues_27; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_28 <= io_adcValues_28; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_29 <= io_adcValues_29; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_30 <= io_adcValues_30; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_31 <= io_adcValues_31; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_32 <= io_adcValues_32; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_33 <= io_adcValues_33; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_34 <= io_adcValues_34; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_35 <= io_adcValues_35; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_36 <= io_adcValues_36; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_37 <= io_adcValues_37; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_38 <= io_adcValues_38; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_39 <= io_adcValues_39; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_40 <= io_adcValues_40; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_41 <= io_adcValues_41; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_42 <= io_adcValues_42; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_43 <= io_adcValues_43; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_44 <= io_adcValues_44; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_45 <= io_adcValues_45; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_46 <= io_adcValues_46; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_47 <= io_adcValues_47; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_48 <= io_adcValues_48; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_49 <= io_adcValues_49; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_50 <= io_adcValues_50; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_51 <= io_adcValues_51; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_52 <= io_adcValues_52; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_53 <= io_adcValues_53; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_54 <= io_adcValues_54; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_55 <= io_adcValues_55; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_56 <= io_adcValues_56; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_57 <= io_adcValues_57; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_58 <= io_adcValues_58; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_59 <= io_adcValues_59; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_60 <= io_adcValues_60; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_61 <= io_adcValues_61; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_62 <= io_adcValues_62; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_63 <= io_adcValues_63; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_64 <= io_adcValues_64; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_65 <= io_adcValues_65; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_66 <= io_adcValues_66; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_67 <= io_adcValues_67; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_68 <= io_adcValues_68; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_69 <= io_adcValues_69; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_70 <= io_adcValues_70; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_71 <= io_adcValues_71; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_72 <= io_adcValues_72; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_73 <= io_adcValues_73; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_74 <= io_adcValues_74; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_75 <= io_adcValues_75; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_76 <= io_adcValues_76; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_77 <= io_adcValues_77; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_78 <= io_adcValues_78; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_79 <= io_adcValues_79; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_80 <= io_adcValues_80; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_81 <= io_adcValues_81; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_82 <= io_adcValues_82; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_83 <= io_adcValues_83; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_84 <= io_adcValues_84; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_85 <= io_adcValues_85; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_86 <= io_adcValues_86; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_87 <= io_adcValues_87; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_88 <= io_adcValues_88; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_89 <= io_adcValues_89; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_90 <= io_adcValues_90; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_91 <= io_adcValues_91; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_92 <= io_adcValues_92; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_93 <= io_adcValues_93; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_94 <= io_adcValues_94; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_95 <= io_adcValues_95; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_96 <= io_adcValues_96; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_97 <= io_adcValues_97; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_98 <= io_adcValues_98; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_99 <= io_adcValues_99; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_100 <= io_adcValues_100; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_101 <= io_adcValues_101; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_102 <= io_adcValues_102; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_103 <= io_adcValues_103; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_104 <= io_adcValues_104; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_105 <= io_adcValues_105; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_106 <= io_adcValues_106; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_107 <= io_adcValues_107; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_108 <= io_adcValues_108; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_109 <= io_adcValues_109; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_110 <= io_adcValues_110; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_111 <= io_adcValues_111; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_112 <= io_adcValues_112; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_113 <= io_adcValues_113; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_114 <= io_adcValues_114; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_115 <= io_adcValues_115; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_116 <= io_adcValues_116; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_117 <= io_adcValues_117; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_118 <= io_adcValues_118; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_119 <= io_adcValues_119; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_120 <= io_adcValues_120; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_121 <= io_adcValues_121; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_122 <= io_adcValues_122; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_123 <= io_adcValues_123; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_124 <= io_adcValues_124; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_125 <= io_adcValues_125; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_126 <= io_adcValues_126; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h4 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_4_127 <= io_adcValues_127; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_0 <= io_adcValues_0; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_1 <= io_adcValues_1; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_2 <= io_adcValues_2; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_3 <= io_adcValues_3; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_4 <= io_adcValues_4; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_5 <= io_adcValues_5; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_6 <= io_adcValues_6; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_7 <= io_adcValues_7; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_8 <= io_adcValues_8; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_9 <= io_adcValues_9; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_10 <= io_adcValues_10; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_11 <= io_adcValues_11; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_12 <= io_adcValues_12; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_13 <= io_adcValues_13; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_14 <= io_adcValues_14; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_15 <= io_adcValues_15; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_16 <= io_adcValues_16; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_17 <= io_adcValues_17; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_18 <= io_adcValues_18; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_19 <= io_adcValues_19; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_20 <= io_adcValues_20; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_21 <= io_adcValues_21; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_22 <= io_adcValues_22; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_23 <= io_adcValues_23; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_24 <= io_adcValues_24; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_25 <= io_adcValues_25; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_26 <= io_adcValues_26; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_27 <= io_adcValues_27; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_28 <= io_adcValues_28; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_29 <= io_adcValues_29; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_30 <= io_adcValues_30; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_31 <= io_adcValues_31; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_32 <= io_adcValues_32; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_33 <= io_adcValues_33; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_34 <= io_adcValues_34; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_35 <= io_adcValues_35; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_36 <= io_adcValues_36; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_37 <= io_adcValues_37; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_38 <= io_adcValues_38; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_39 <= io_adcValues_39; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_40 <= io_adcValues_40; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_41 <= io_adcValues_41; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_42 <= io_adcValues_42; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_43 <= io_adcValues_43; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_44 <= io_adcValues_44; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_45 <= io_adcValues_45; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_46 <= io_adcValues_46; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_47 <= io_adcValues_47; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_48 <= io_adcValues_48; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_49 <= io_adcValues_49; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_50 <= io_adcValues_50; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_51 <= io_adcValues_51; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_52 <= io_adcValues_52; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_53 <= io_adcValues_53; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_54 <= io_adcValues_54; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_55 <= io_adcValues_55; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_56 <= io_adcValues_56; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_57 <= io_adcValues_57; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_58 <= io_adcValues_58; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_59 <= io_adcValues_59; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_60 <= io_adcValues_60; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_61 <= io_adcValues_61; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_62 <= io_adcValues_62; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_63 <= io_adcValues_63; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_64 <= io_adcValues_64; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_65 <= io_adcValues_65; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_66 <= io_adcValues_66; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_67 <= io_adcValues_67; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_68 <= io_adcValues_68; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_69 <= io_adcValues_69; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_70 <= io_adcValues_70; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_71 <= io_adcValues_71; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_72 <= io_adcValues_72; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_73 <= io_adcValues_73; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_74 <= io_adcValues_74; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_75 <= io_adcValues_75; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_76 <= io_adcValues_76; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_77 <= io_adcValues_77; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_78 <= io_adcValues_78; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_79 <= io_adcValues_79; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_80 <= io_adcValues_80; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_81 <= io_adcValues_81; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_82 <= io_adcValues_82; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_83 <= io_adcValues_83; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_84 <= io_adcValues_84; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_85 <= io_adcValues_85; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_86 <= io_adcValues_86; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_87 <= io_adcValues_87; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_88 <= io_adcValues_88; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_89 <= io_adcValues_89; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_90 <= io_adcValues_90; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_91 <= io_adcValues_91; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_92 <= io_adcValues_92; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_93 <= io_adcValues_93; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_94 <= io_adcValues_94; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_95 <= io_adcValues_95; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_96 <= io_adcValues_96; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_97 <= io_adcValues_97; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_98 <= io_adcValues_98; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_99 <= io_adcValues_99; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_100 <= io_adcValues_100; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_101 <= io_adcValues_101; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_102 <= io_adcValues_102; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_103 <= io_adcValues_103; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_104 <= io_adcValues_104; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_105 <= io_adcValues_105; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_106 <= io_adcValues_106; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_107 <= io_adcValues_107; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_108 <= io_adcValues_108; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_109 <= io_adcValues_109; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_110 <= io_adcValues_110; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_111 <= io_adcValues_111; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_112 <= io_adcValues_112; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_113 <= io_adcValues_113; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_114 <= io_adcValues_114; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_115 <= io_adcValues_115; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_116 <= io_adcValues_116; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_117 <= io_adcValues_117; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_118 <= io_adcValues_118; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_119 <= io_adcValues_119; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_120 <= io_adcValues_120; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_121 <= io_adcValues_121; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_122 <= io_adcValues_122; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_123 <= io_adcValues_123; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_124 <= io_adcValues_124; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_125 <= io_adcValues_125; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_126 <= io_adcValues_126; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h5 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_5_127 <= io_adcValues_127; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_0 <= io_adcValues_0; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_1 <= io_adcValues_1; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_2 <= io_adcValues_2; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_3 <= io_adcValues_3; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_4 <= io_adcValues_4; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_5 <= io_adcValues_5; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_6 <= io_adcValues_6; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_7 <= io_adcValues_7; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_8 <= io_adcValues_8; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_9 <= io_adcValues_9; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_10 <= io_adcValues_10; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_11 <= io_adcValues_11; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_12 <= io_adcValues_12; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_13 <= io_adcValues_13; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_14 <= io_adcValues_14; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_15 <= io_adcValues_15; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_16 <= io_adcValues_16; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_17 <= io_adcValues_17; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_18 <= io_adcValues_18; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_19 <= io_adcValues_19; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_20 <= io_adcValues_20; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_21 <= io_adcValues_21; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_22 <= io_adcValues_22; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_23 <= io_adcValues_23; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_24 <= io_adcValues_24; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_25 <= io_adcValues_25; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_26 <= io_adcValues_26; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_27 <= io_adcValues_27; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_28 <= io_adcValues_28; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_29 <= io_adcValues_29; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_30 <= io_adcValues_30; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_31 <= io_adcValues_31; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_32 <= io_adcValues_32; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_33 <= io_adcValues_33; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_34 <= io_adcValues_34; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_35 <= io_adcValues_35; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_36 <= io_adcValues_36; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_37 <= io_adcValues_37; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_38 <= io_adcValues_38; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_39 <= io_adcValues_39; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_40 <= io_adcValues_40; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_41 <= io_adcValues_41; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_42 <= io_adcValues_42; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_43 <= io_adcValues_43; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_44 <= io_adcValues_44; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_45 <= io_adcValues_45; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_46 <= io_adcValues_46; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_47 <= io_adcValues_47; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_48 <= io_adcValues_48; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_49 <= io_adcValues_49; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_50 <= io_adcValues_50; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_51 <= io_adcValues_51; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_52 <= io_adcValues_52; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_53 <= io_adcValues_53; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_54 <= io_adcValues_54; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_55 <= io_adcValues_55; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_56 <= io_adcValues_56; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_57 <= io_adcValues_57; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_58 <= io_adcValues_58; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_59 <= io_adcValues_59; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_60 <= io_adcValues_60; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_61 <= io_adcValues_61; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_62 <= io_adcValues_62; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_63 <= io_adcValues_63; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_64 <= io_adcValues_64; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_65 <= io_adcValues_65; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_66 <= io_adcValues_66; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_67 <= io_adcValues_67; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_68 <= io_adcValues_68; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_69 <= io_adcValues_69; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_70 <= io_adcValues_70; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_71 <= io_adcValues_71; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_72 <= io_adcValues_72; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_73 <= io_adcValues_73; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_74 <= io_adcValues_74; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_75 <= io_adcValues_75; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_76 <= io_adcValues_76; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_77 <= io_adcValues_77; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_78 <= io_adcValues_78; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_79 <= io_adcValues_79; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_80 <= io_adcValues_80; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_81 <= io_adcValues_81; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_82 <= io_adcValues_82; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_83 <= io_adcValues_83; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_84 <= io_adcValues_84; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_85 <= io_adcValues_85; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_86 <= io_adcValues_86; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_87 <= io_adcValues_87; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_88 <= io_adcValues_88; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_89 <= io_adcValues_89; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_90 <= io_adcValues_90; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_91 <= io_adcValues_91; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_92 <= io_adcValues_92; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_93 <= io_adcValues_93; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_94 <= io_adcValues_94; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_95 <= io_adcValues_95; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_96 <= io_adcValues_96; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_97 <= io_adcValues_97; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_98 <= io_adcValues_98; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_99 <= io_adcValues_99; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_100 <= io_adcValues_100; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_101 <= io_adcValues_101; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_102 <= io_adcValues_102; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_103 <= io_adcValues_103; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_104 <= io_adcValues_104; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_105 <= io_adcValues_105; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_106 <= io_adcValues_106; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_107 <= io_adcValues_107; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_108 <= io_adcValues_108; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_109 <= io_adcValues_109; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_110 <= io_adcValues_110; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_111 <= io_adcValues_111; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_112 <= io_adcValues_112; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_113 <= io_adcValues_113; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_114 <= io_adcValues_114; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_115 <= io_adcValues_115; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_116 <= io_adcValues_116; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_117 <= io_adcValues_117; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_118 <= io_adcValues_118; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_119 <= io_adcValues_119; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_120 <= io_adcValues_120; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_121 <= io_adcValues_121; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_122 <= io_adcValues_122; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_123 <= io_adcValues_123; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_124 <= io_adcValues_124; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_125 <= io_adcValues_125; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_126 <= io_adcValues_126; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h6 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_6_127 <= io_adcValues_127; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_0 <= io_adcValues_0; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_1 <= io_adcValues_1; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_2 <= io_adcValues_2; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_3 <= io_adcValues_3; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_4 <= io_adcValues_4; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_5 <= io_adcValues_5; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_6 <= io_adcValues_6; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_7 <= io_adcValues_7; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_8 <= io_adcValues_8; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_9 <= io_adcValues_9; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_10 <= io_adcValues_10; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_11 <= io_adcValues_11; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_12 <= io_adcValues_12; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_13 <= io_adcValues_13; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_14 <= io_adcValues_14; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_15 <= io_adcValues_15; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_16 <= io_adcValues_16; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_17 <= io_adcValues_17; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_18 <= io_adcValues_18; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_19 <= io_adcValues_19; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_20 <= io_adcValues_20; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_21 <= io_adcValues_21; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_22 <= io_adcValues_22; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_23 <= io_adcValues_23; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_24 <= io_adcValues_24; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_25 <= io_adcValues_25; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_26 <= io_adcValues_26; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_27 <= io_adcValues_27; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_28 <= io_adcValues_28; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_29 <= io_adcValues_29; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_30 <= io_adcValues_30; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_31 <= io_adcValues_31; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_32 <= io_adcValues_32; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_33 <= io_adcValues_33; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_34 <= io_adcValues_34; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_35 <= io_adcValues_35; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_36 <= io_adcValues_36; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_37 <= io_adcValues_37; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_38 <= io_adcValues_38; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_39 <= io_adcValues_39; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_40 <= io_adcValues_40; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_41 <= io_adcValues_41; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_42 <= io_adcValues_42; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_43 <= io_adcValues_43; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_44 <= io_adcValues_44; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_45 <= io_adcValues_45; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_46 <= io_adcValues_46; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_47 <= io_adcValues_47; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_48 <= io_adcValues_48; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_49 <= io_adcValues_49; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_50 <= io_adcValues_50; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_51 <= io_adcValues_51; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_52 <= io_adcValues_52; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_53 <= io_adcValues_53; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_54 <= io_adcValues_54; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_55 <= io_adcValues_55; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_56 <= io_adcValues_56; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_57 <= io_adcValues_57; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_58 <= io_adcValues_58; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_59 <= io_adcValues_59; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_60 <= io_adcValues_60; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_61 <= io_adcValues_61; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_62 <= io_adcValues_62; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_63 <= io_adcValues_63; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_64 <= io_adcValues_64; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_65 <= io_adcValues_65; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_66 <= io_adcValues_66; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_67 <= io_adcValues_67; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_68 <= io_adcValues_68; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_69 <= io_adcValues_69; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_70 <= io_adcValues_70; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_71 <= io_adcValues_71; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_72 <= io_adcValues_72; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_73 <= io_adcValues_73; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_74 <= io_adcValues_74; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_75 <= io_adcValues_75; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_76 <= io_adcValues_76; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_77 <= io_adcValues_77; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_78 <= io_adcValues_78; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_79 <= io_adcValues_79; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_80 <= io_adcValues_80; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_81 <= io_adcValues_81; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_82 <= io_adcValues_82; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_83 <= io_adcValues_83; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_84 <= io_adcValues_84; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_85 <= io_adcValues_85; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_86 <= io_adcValues_86; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_87 <= io_adcValues_87; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_88 <= io_adcValues_88; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_89 <= io_adcValues_89; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_90 <= io_adcValues_90; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_91 <= io_adcValues_91; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_92 <= io_adcValues_92; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_93 <= io_adcValues_93; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_94 <= io_adcValues_94; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_95 <= io_adcValues_95; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_96 <= io_adcValues_96; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_97 <= io_adcValues_97; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_98 <= io_adcValues_98; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_99 <= io_adcValues_99; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_100 <= io_adcValues_100; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_101 <= io_adcValues_101; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_102 <= io_adcValues_102; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_103 <= io_adcValues_103; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_104 <= io_adcValues_104; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_105 <= io_adcValues_105; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_106 <= io_adcValues_106; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_107 <= io_adcValues_107; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_108 <= io_adcValues_108; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_109 <= io_adcValues_109; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_110 <= io_adcValues_110; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_111 <= io_adcValues_111; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_112 <= io_adcValues_112; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_113 <= io_adcValues_113; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_114 <= io_adcValues_114; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_115 <= io_adcValues_115; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_116 <= io_adcValues_116; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_117 <= io_adcValues_117; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_118 <= io_adcValues_118; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_119 <= io_adcValues_119; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_120 <= io_adcValues_120; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_121 <= io_adcValues_121; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_122 <= io_adcValues_122; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_123 <= io_adcValues_123; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_124 <= io_adcValues_124; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_125 <= io_adcValues_125; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_126 <= io_adcValues_126; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h7 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_7_127 <= io_adcValues_127; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_0 <= io_adcValues_0; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_1 <= io_adcValues_1; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_2 <= io_adcValues_2; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_3 <= io_adcValues_3; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_4 <= io_adcValues_4; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_5 <= io_adcValues_5; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_6 <= io_adcValues_6; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_7 <= io_adcValues_7; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_8 <= io_adcValues_8; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_9 <= io_adcValues_9; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_10 <= io_adcValues_10; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_11 <= io_adcValues_11; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_12 <= io_adcValues_12; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_13 <= io_adcValues_13; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_14 <= io_adcValues_14; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_15 <= io_adcValues_15; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_16 <= io_adcValues_16; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_17 <= io_adcValues_17; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_18 <= io_adcValues_18; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_19 <= io_adcValues_19; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_20 <= io_adcValues_20; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_21 <= io_adcValues_21; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_22 <= io_adcValues_22; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_23 <= io_adcValues_23; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_24 <= io_adcValues_24; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_25 <= io_adcValues_25; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_26 <= io_adcValues_26; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_27 <= io_adcValues_27; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_28 <= io_adcValues_28; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_29 <= io_adcValues_29; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_30 <= io_adcValues_30; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_31 <= io_adcValues_31; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_32 <= io_adcValues_32; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_33 <= io_adcValues_33; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_34 <= io_adcValues_34; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_35 <= io_adcValues_35; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_36 <= io_adcValues_36; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_37 <= io_adcValues_37; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_38 <= io_adcValues_38; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_39 <= io_adcValues_39; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_40 <= io_adcValues_40; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_41 <= io_adcValues_41; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_42 <= io_adcValues_42; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_43 <= io_adcValues_43; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_44 <= io_adcValues_44; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_45 <= io_adcValues_45; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_46 <= io_adcValues_46; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_47 <= io_adcValues_47; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_48 <= io_adcValues_48; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_49 <= io_adcValues_49; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_50 <= io_adcValues_50; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_51 <= io_adcValues_51; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_52 <= io_adcValues_52; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_53 <= io_adcValues_53; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_54 <= io_adcValues_54; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_55 <= io_adcValues_55; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_56 <= io_adcValues_56; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_57 <= io_adcValues_57; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_58 <= io_adcValues_58; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_59 <= io_adcValues_59; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_60 <= io_adcValues_60; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_61 <= io_adcValues_61; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_62 <= io_adcValues_62; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_63 <= io_adcValues_63; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_64 <= io_adcValues_64; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_65 <= io_adcValues_65; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_66 <= io_adcValues_66; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_67 <= io_adcValues_67; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_68 <= io_adcValues_68; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_69 <= io_adcValues_69; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_70 <= io_adcValues_70; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_71 <= io_adcValues_71; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_72 <= io_adcValues_72; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_73 <= io_adcValues_73; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_74 <= io_adcValues_74; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_75 <= io_adcValues_75; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_76 <= io_adcValues_76; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_77 <= io_adcValues_77; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_78 <= io_adcValues_78; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_79 <= io_adcValues_79; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_80 <= io_adcValues_80; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_81 <= io_adcValues_81; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_82 <= io_adcValues_82; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_83 <= io_adcValues_83; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_84 <= io_adcValues_84; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_85 <= io_adcValues_85; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_86 <= io_adcValues_86; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_87 <= io_adcValues_87; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_88 <= io_adcValues_88; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_89 <= io_adcValues_89; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_90 <= io_adcValues_90; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_91 <= io_adcValues_91; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_92 <= io_adcValues_92; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_93 <= io_adcValues_93; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_94 <= io_adcValues_94; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_95 <= io_adcValues_95; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_96 <= io_adcValues_96; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_97 <= io_adcValues_97; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_98 <= io_adcValues_98; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_99 <= io_adcValues_99; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_100 <= io_adcValues_100; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_101 <= io_adcValues_101; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_102 <= io_adcValues_102; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_103 <= io_adcValues_103; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_104 <= io_adcValues_104; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_105 <= io_adcValues_105; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_106 <= io_adcValues_106; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_107 <= io_adcValues_107; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_108 <= io_adcValues_108; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_109 <= io_adcValues_109; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_110 <= io_adcValues_110; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_111 <= io_adcValues_111; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_112 <= io_adcValues_112; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_113 <= io_adcValues_113; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_114 <= io_adcValues_114; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_115 <= io_adcValues_115; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_116 <= io_adcValues_116; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_117 <= io_adcValues_117; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_118 <= io_adcValues_118; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_119 <= io_adcValues_119; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_120 <= io_adcValues_120; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_121 <= io_adcValues_121; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_122 <= io_adcValues_122; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_123 <= io_adcValues_123; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_124 <= io_adcValues_124; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_125 <= io_adcValues_125; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_126 <= io_adcValues_126; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h8 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_8_127 <= io_adcValues_127; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_0 <= io_adcValues_0; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_1 <= io_adcValues_1; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_2 <= io_adcValues_2; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_3 <= io_adcValues_3; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_4 <= io_adcValues_4; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_5 <= io_adcValues_5; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_6 <= io_adcValues_6; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_7 <= io_adcValues_7; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_8 <= io_adcValues_8; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_9 <= io_adcValues_9; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_10 <= io_adcValues_10; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_11 <= io_adcValues_11; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_12 <= io_adcValues_12; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_13 <= io_adcValues_13; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_14 <= io_adcValues_14; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_15 <= io_adcValues_15; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_16 <= io_adcValues_16; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_17 <= io_adcValues_17; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_18 <= io_adcValues_18; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_19 <= io_adcValues_19; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_20 <= io_adcValues_20; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_21 <= io_adcValues_21; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_22 <= io_adcValues_22; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_23 <= io_adcValues_23; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_24 <= io_adcValues_24; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_25 <= io_adcValues_25; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_26 <= io_adcValues_26; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_27 <= io_adcValues_27; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_28 <= io_adcValues_28; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_29 <= io_adcValues_29; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_30 <= io_adcValues_30; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_31 <= io_adcValues_31; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_32 <= io_adcValues_32; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_33 <= io_adcValues_33; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_34 <= io_adcValues_34; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_35 <= io_adcValues_35; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_36 <= io_adcValues_36; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_37 <= io_adcValues_37; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_38 <= io_adcValues_38; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_39 <= io_adcValues_39; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_40 <= io_adcValues_40; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_41 <= io_adcValues_41; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_42 <= io_adcValues_42; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_43 <= io_adcValues_43; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_44 <= io_adcValues_44; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_45 <= io_adcValues_45; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_46 <= io_adcValues_46; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_47 <= io_adcValues_47; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_48 <= io_adcValues_48; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_49 <= io_adcValues_49; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_50 <= io_adcValues_50; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_51 <= io_adcValues_51; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_52 <= io_adcValues_52; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_53 <= io_adcValues_53; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_54 <= io_adcValues_54; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_55 <= io_adcValues_55; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_56 <= io_adcValues_56; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_57 <= io_adcValues_57; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_58 <= io_adcValues_58; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_59 <= io_adcValues_59; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_60 <= io_adcValues_60; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_61 <= io_adcValues_61; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_62 <= io_adcValues_62; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_63 <= io_adcValues_63; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_64 <= io_adcValues_64; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_65 <= io_adcValues_65; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_66 <= io_adcValues_66; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_67 <= io_adcValues_67; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_68 <= io_adcValues_68; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_69 <= io_adcValues_69; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_70 <= io_adcValues_70; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_71 <= io_adcValues_71; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_72 <= io_adcValues_72; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_73 <= io_adcValues_73; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_74 <= io_adcValues_74; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_75 <= io_adcValues_75; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_76 <= io_adcValues_76; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_77 <= io_adcValues_77; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_78 <= io_adcValues_78; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_79 <= io_adcValues_79; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_80 <= io_adcValues_80; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_81 <= io_adcValues_81; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_82 <= io_adcValues_82; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_83 <= io_adcValues_83; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_84 <= io_adcValues_84; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_85 <= io_adcValues_85; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_86 <= io_adcValues_86; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_87 <= io_adcValues_87; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_88 <= io_adcValues_88; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_89 <= io_adcValues_89; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_90 <= io_adcValues_90; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_91 <= io_adcValues_91; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_92 <= io_adcValues_92; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_93 <= io_adcValues_93; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_94 <= io_adcValues_94; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_95 <= io_adcValues_95; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_96 <= io_adcValues_96; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_97 <= io_adcValues_97; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_98 <= io_adcValues_98; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_99 <= io_adcValues_99; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_100 <= io_adcValues_100; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_101 <= io_adcValues_101; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_102 <= io_adcValues_102; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_103 <= io_adcValues_103; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_104 <= io_adcValues_104; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_105 <= io_adcValues_105; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_106 <= io_adcValues_106; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_107 <= io_adcValues_107; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_108 <= io_adcValues_108; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_109 <= io_adcValues_109; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_110 <= io_adcValues_110; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_111 <= io_adcValues_111; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_112 <= io_adcValues_112; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_113 <= io_adcValues_113; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_114 <= io_adcValues_114; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_115 <= io_adcValues_115; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_116 <= io_adcValues_116; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_117 <= io_adcValues_117; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_118 <= io_adcValues_118; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_119 <= io_adcValues_119; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_120 <= io_adcValues_120; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_121 <= io_adcValues_121; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_122 <= io_adcValues_122; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_123 <= io_adcValues_123; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_124 <= io_adcValues_124; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_125 <= io_adcValues_125; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_126 <= io_adcValues_126; // @[BufferAMSNew.scala 24:28]
    end
    if (4'h9 == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_9_127 <= io_adcValues_127; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_0 <= io_adcValues_0; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_1 <= io_adcValues_1; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_2 <= io_adcValues_2; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_3 <= io_adcValues_3; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_4 <= io_adcValues_4; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_5 <= io_adcValues_5; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_6 <= io_adcValues_6; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_7 <= io_adcValues_7; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_8 <= io_adcValues_8; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_9 <= io_adcValues_9; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_10 <= io_adcValues_10; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_11 <= io_adcValues_11; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_12 <= io_adcValues_12; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_13 <= io_adcValues_13; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_14 <= io_adcValues_14; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_15 <= io_adcValues_15; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_16 <= io_adcValues_16; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_17 <= io_adcValues_17; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_18 <= io_adcValues_18; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_19 <= io_adcValues_19; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_20 <= io_adcValues_20; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_21 <= io_adcValues_21; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_22 <= io_adcValues_22; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_23 <= io_adcValues_23; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_24 <= io_adcValues_24; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_25 <= io_adcValues_25; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_26 <= io_adcValues_26; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_27 <= io_adcValues_27; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_28 <= io_adcValues_28; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_29 <= io_adcValues_29; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_30 <= io_adcValues_30; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_31 <= io_adcValues_31; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_32 <= io_adcValues_32; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_33 <= io_adcValues_33; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_34 <= io_adcValues_34; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_35 <= io_adcValues_35; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_36 <= io_adcValues_36; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_37 <= io_adcValues_37; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_38 <= io_adcValues_38; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_39 <= io_adcValues_39; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_40 <= io_adcValues_40; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_41 <= io_adcValues_41; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_42 <= io_adcValues_42; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_43 <= io_adcValues_43; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_44 <= io_adcValues_44; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_45 <= io_adcValues_45; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_46 <= io_adcValues_46; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_47 <= io_adcValues_47; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_48 <= io_adcValues_48; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_49 <= io_adcValues_49; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_50 <= io_adcValues_50; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_51 <= io_adcValues_51; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_52 <= io_adcValues_52; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_53 <= io_adcValues_53; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_54 <= io_adcValues_54; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_55 <= io_adcValues_55; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_56 <= io_adcValues_56; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_57 <= io_adcValues_57; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_58 <= io_adcValues_58; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_59 <= io_adcValues_59; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_60 <= io_adcValues_60; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_61 <= io_adcValues_61; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_62 <= io_adcValues_62; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_63 <= io_adcValues_63; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_64 <= io_adcValues_64; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_65 <= io_adcValues_65; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_66 <= io_adcValues_66; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_67 <= io_adcValues_67; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_68 <= io_adcValues_68; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_69 <= io_adcValues_69; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_70 <= io_adcValues_70; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_71 <= io_adcValues_71; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_72 <= io_adcValues_72; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_73 <= io_adcValues_73; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_74 <= io_adcValues_74; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_75 <= io_adcValues_75; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_76 <= io_adcValues_76; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_77 <= io_adcValues_77; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_78 <= io_adcValues_78; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_79 <= io_adcValues_79; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_80 <= io_adcValues_80; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_81 <= io_adcValues_81; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_82 <= io_adcValues_82; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_83 <= io_adcValues_83; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_84 <= io_adcValues_84; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_85 <= io_adcValues_85; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_86 <= io_adcValues_86; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_87 <= io_adcValues_87; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_88 <= io_adcValues_88; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_89 <= io_adcValues_89; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_90 <= io_adcValues_90; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_91 <= io_adcValues_91; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_92 <= io_adcValues_92; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_93 <= io_adcValues_93; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_94 <= io_adcValues_94; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_95 <= io_adcValues_95; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_96 <= io_adcValues_96; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_97 <= io_adcValues_97; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_98 <= io_adcValues_98; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_99 <= io_adcValues_99; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_100 <= io_adcValues_100; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_101 <= io_adcValues_101; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_102 <= io_adcValues_102; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_103 <= io_adcValues_103; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_104 <= io_adcValues_104; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_105 <= io_adcValues_105; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_106 <= io_adcValues_106; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_107 <= io_adcValues_107; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_108 <= io_adcValues_108; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_109 <= io_adcValues_109; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_110 <= io_adcValues_110; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_111 <= io_adcValues_111; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_112 <= io_adcValues_112; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_113 <= io_adcValues_113; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_114 <= io_adcValues_114; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_115 <= io_adcValues_115; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_116 <= io_adcValues_116; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_117 <= io_adcValues_117; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_118 <= io_adcValues_118; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_119 <= io_adcValues_119; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_120 <= io_adcValues_120; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_121 <= io_adcValues_121; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_122 <= io_adcValues_122; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_123 <= io_adcValues_123; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_124 <= io_adcValues_124; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_125 <= io_adcValues_125; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_126 <= io_adcValues_126; // @[BufferAMSNew.scala 24:28]
    end
    if (4'ha == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_10_127 <= io_adcValues_127; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_0 <= io_adcValues_0; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_1 <= io_adcValues_1; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_2 <= io_adcValues_2; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_3 <= io_adcValues_3; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_4 <= io_adcValues_4; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_5 <= io_adcValues_5; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_6 <= io_adcValues_6; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_7 <= io_adcValues_7; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_8 <= io_adcValues_8; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_9 <= io_adcValues_9; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_10 <= io_adcValues_10; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_11 <= io_adcValues_11; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_12 <= io_adcValues_12; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_13 <= io_adcValues_13; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_14 <= io_adcValues_14; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_15 <= io_adcValues_15; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_16 <= io_adcValues_16; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_17 <= io_adcValues_17; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_18 <= io_adcValues_18; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_19 <= io_adcValues_19; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_20 <= io_adcValues_20; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_21 <= io_adcValues_21; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_22 <= io_adcValues_22; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_23 <= io_adcValues_23; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_24 <= io_adcValues_24; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_25 <= io_adcValues_25; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_26 <= io_adcValues_26; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_27 <= io_adcValues_27; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_28 <= io_adcValues_28; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_29 <= io_adcValues_29; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_30 <= io_adcValues_30; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_31 <= io_adcValues_31; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_32 <= io_adcValues_32; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_33 <= io_adcValues_33; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_34 <= io_adcValues_34; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_35 <= io_adcValues_35; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_36 <= io_adcValues_36; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_37 <= io_adcValues_37; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_38 <= io_adcValues_38; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_39 <= io_adcValues_39; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_40 <= io_adcValues_40; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_41 <= io_adcValues_41; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_42 <= io_adcValues_42; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_43 <= io_adcValues_43; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_44 <= io_adcValues_44; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_45 <= io_adcValues_45; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_46 <= io_adcValues_46; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_47 <= io_adcValues_47; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_48 <= io_adcValues_48; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_49 <= io_adcValues_49; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_50 <= io_adcValues_50; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_51 <= io_adcValues_51; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_52 <= io_adcValues_52; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_53 <= io_adcValues_53; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_54 <= io_adcValues_54; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_55 <= io_adcValues_55; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_56 <= io_adcValues_56; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_57 <= io_adcValues_57; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_58 <= io_adcValues_58; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_59 <= io_adcValues_59; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_60 <= io_adcValues_60; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_61 <= io_adcValues_61; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_62 <= io_adcValues_62; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_63 <= io_adcValues_63; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_64 <= io_adcValues_64; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_65 <= io_adcValues_65; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_66 <= io_adcValues_66; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_67 <= io_adcValues_67; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_68 <= io_adcValues_68; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_69 <= io_adcValues_69; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_70 <= io_adcValues_70; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_71 <= io_adcValues_71; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_72 <= io_adcValues_72; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_73 <= io_adcValues_73; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_74 <= io_adcValues_74; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_75 <= io_adcValues_75; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_76 <= io_adcValues_76; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_77 <= io_adcValues_77; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_78 <= io_adcValues_78; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_79 <= io_adcValues_79; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_80 <= io_adcValues_80; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_81 <= io_adcValues_81; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_82 <= io_adcValues_82; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_83 <= io_adcValues_83; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_84 <= io_adcValues_84; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_85 <= io_adcValues_85; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_86 <= io_adcValues_86; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_87 <= io_adcValues_87; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_88 <= io_adcValues_88; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_89 <= io_adcValues_89; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_90 <= io_adcValues_90; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_91 <= io_adcValues_91; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_92 <= io_adcValues_92; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_93 <= io_adcValues_93; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_94 <= io_adcValues_94; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_95 <= io_adcValues_95; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_96 <= io_adcValues_96; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_97 <= io_adcValues_97; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_98 <= io_adcValues_98; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_99 <= io_adcValues_99; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_100 <= io_adcValues_100; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_101 <= io_adcValues_101; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_102 <= io_adcValues_102; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_103 <= io_adcValues_103; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_104 <= io_adcValues_104; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_105 <= io_adcValues_105; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_106 <= io_adcValues_106; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_107 <= io_adcValues_107; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_108 <= io_adcValues_108; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_109 <= io_adcValues_109; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_110 <= io_adcValues_110; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_111 <= io_adcValues_111; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_112 <= io_adcValues_112; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_113 <= io_adcValues_113; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_114 <= io_adcValues_114; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_115 <= io_adcValues_115; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_116 <= io_adcValues_116; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_117 <= io_adcValues_117; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_118 <= io_adcValues_118; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_119 <= io_adcValues_119; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_120 <= io_adcValues_120; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_121 <= io_adcValues_121; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_122 <= io_adcValues_122; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_123 <= io_adcValues_123; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_124 <= io_adcValues_124; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_125 <= io_adcValues_125; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_126 <= io_adcValues_126; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hb == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_11_127 <= io_adcValues_127; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_0 <= io_adcValues_0; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_1 <= io_adcValues_1; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_2 <= io_adcValues_2; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_3 <= io_adcValues_3; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_4 <= io_adcValues_4; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_5 <= io_adcValues_5; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_6 <= io_adcValues_6; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_7 <= io_adcValues_7; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_8 <= io_adcValues_8; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_9 <= io_adcValues_9; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_10 <= io_adcValues_10; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_11 <= io_adcValues_11; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_12 <= io_adcValues_12; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_13 <= io_adcValues_13; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_14 <= io_adcValues_14; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_15 <= io_adcValues_15; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_16 <= io_adcValues_16; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_17 <= io_adcValues_17; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_18 <= io_adcValues_18; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_19 <= io_adcValues_19; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_20 <= io_adcValues_20; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_21 <= io_adcValues_21; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_22 <= io_adcValues_22; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_23 <= io_adcValues_23; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_24 <= io_adcValues_24; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_25 <= io_adcValues_25; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_26 <= io_adcValues_26; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_27 <= io_adcValues_27; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_28 <= io_adcValues_28; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_29 <= io_adcValues_29; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_30 <= io_adcValues_30; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_31 <= io_adcValues_31; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_32 <= io_adcValues_32; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_33 <= io_adcValues_33; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_34 <= io_adcValues_34; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_35 <= io_adcValues_35; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_36 <= io_adcValues_36; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_37 <= io_adcValues_37; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_38 <= io_adcValues_38; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_39 <= io_adcValues_39; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_40 <= io_adcValues_40; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_41 <= io_adcValues_41; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_42 <= io_adcValues_42; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_43 <= io_adcValues_43; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_44 <= io_adcValues_44; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_45 <= io_adcValues_45; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_46 <= io_adcValues_46; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_47 <= io_adcValues_47; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_48 <= io_adcValues_48; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_49 <= io_adcValues_49; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_50 <= io_adcValues_50; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_51 <= io_adcValues_51; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_52 <= io_adcValues_52; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_53 <= io_adcValues_53; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_54 <= io_adcValues_54; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_55 <= io_adcValues_55; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_56 <= io_adcValues_56; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_57 <= io_adcValues_57; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_58 <= io_adcValues_58; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_59 <= io_adcValues_59; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_60 <= io_adcValues_60; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_61 <= io_adcValues_61; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_62 <= io_adcValues_62; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_63 <= io_adcValues_63; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_64 <= io_adcValues_64; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_65 <= io_adcValues_65; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_66 <= io_adcValues_66; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_67 <= io_adcValues_67; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_68 <= io_adcValues_68; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_69 <= io_adcValues_69; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_70 <= io_adcValues_70; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_71 <= io_adcValues_71; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_72 <= io_adcValues_72; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_73 <= io_adcValues_73; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_74 <= io_adcValues_74; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_75 <= io_adcValues_75; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_76 <= io_adcValues_76; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_77 <= io_adcValues_77; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_78 <= io_adcValues_78; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_79 <= io_adcValues_79; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_80 <= io_adcValues_80; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_81 <= io_adcValues_81; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_82 <= io_adcValues_82; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_83 <= io_adcValues_83; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_84 <= io_adcValues_84; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_85 <= io_adcValues_85; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_86 <= io_adcValues_86; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_87 <= io_adcValues_87; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_88 <= io_adcValues_88; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_89 <= io_adcValues_89; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_90 <= io_adcValues_90; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_91 <= io_adcValues_91; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_92 <= io_adcValues_92; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_93 <= io_adcValues_93; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_94 <= io_adcValues_94; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_95 <= io_adcValues_95; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_96 <= io_adcValues_96; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_97 <= io_adcValues_97; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_98 <= io_adcValues_98; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_99 <= io_adcValues_99; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_100 <= io_adcValues_100; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_101 <= io_adcValues_101; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_102 <= io_adcValues_102; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_103 <= io_adcValues_103; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_104 <= io_adcValues_104; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_105 <= io_adcValues_105; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_106 <= io_adcValues_106; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_107 <= io_adcValues_107; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_108 <= io_adcValues_108; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_109 <= io_adcValues_109; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_110 <= io_adcValues_110; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_111 <= io_adcValues_111; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_112 <= io_adcValues_112; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_113 <= io_adcValues_113; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_114 <= io_adcValues_114; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_115 <= io_adcValues_115; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_116 <= io_adcValues_116; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_117 <= io_adcValues_117; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_118 <= io_adcValues_118; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_119 <= io_adcValues_119; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_120 <= io_adcValues_120; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_121 <= io_adcValues_121; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_122 <= io_adcValues_122; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_123 <= io_adcValues_123; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_124 <= io_adcValues_124; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_125 <= io_adcValues_125; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_126 <= io_adcValues_126; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hc == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_12_127 <= io_adcValues_127; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_0 <= io_adcValues_0; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_1 <= io_adcValues_1; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_2 <= io_adcValues_2; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_3 <= io_adcValues_3; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_4 <= io_adcValues_4; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_5 <= io_adcValues_5; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_6 <= io_adcValues_6; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_7 <= io_adcValues_7; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_8 <= io_adcValues_8; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_9 <= io_adcValues_9; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_10 <= io_adcValues_10; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_11 <= io_adcValues_11; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_12 <= io_adcValues_12; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_13 <= io_adcValues_13; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_14 <= io_adcValues_14; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_15 <= io_adcValues_15; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_16 <= io_adcValues_16; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_17 <= io_adcValues_17; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_18 <= io_adcValues_18; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_19 <= io_adcValues_19; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_20 <= io_adcValues_20; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_21 <= io_adcValues_21; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_22 <= io_adcValues_22; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_23 <= io_adcValues_23; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_24 <= io_adcValues_24; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_25 <= io_adcValues_25; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_26 <= io_adcValues_26; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_27 <= io_adcValues_27; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_28 <= io_adcValues_28; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_29 <= io_adcValues_29; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_30 <= io_adcValues_30; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_31 <= io_adcValues_31; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_32 <= io_adcValues_32; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_33 <= io_adcValues_33; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_34 <= io_adcValues_34; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_35 <= io_adcValues_35; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_36 <= io_adcValues_36; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_37 <= io_adcValues_37; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_38 <= io_adcValues_38; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_39 <= io_adcValues_39; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_40 <= io_adcValues_40; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_41 <= io_adcValues_41; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_42 <= io_adcValues_42; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_43 <= io_adcValues_43; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_44 <= io_adcValues_44; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_45 <= io_adcValues_45; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_46 <= io_adcValues_46; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_47 <= io_adcValues_47; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_48 <= io_adcValues_48; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_49 <= io_adcValues_49; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_50 <= io_adcValues_50; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_51 <= io_adcValues_51; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_52 <= io_adcValues_52; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_53 <= io_adcValues_53; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_54 <= io_adcValues_54; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_55 <= io_adcValues_55; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_56 <= io_adcValues_56; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_57 <= io_adcValues_57; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_58 <= io_adcValues_58; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_59 <= io_adcValues_59; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_60 <= io_adcValues_60; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_61 <= io_adcValues_61; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_62 <= io_adcValues_62; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_63 <= io_adcValues_63; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_64 <= io_adcValues_64; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_65 <= io_adcValues_65; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_66 <= io_adcValues_66; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_67 <= io_adcValues_67; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_68 <= io_adcValues_68; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_69 <= io_adcValues_69; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_70 <= io_adcValues_70; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_71 <= io_adcValues_71; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_72 <= io_adcValues_72; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_73 <= io_adcValues_73; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_74 <= io_adcValues_74; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_75 <= io_adcValues_75; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_76 <= io_adcValues_76; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_77 <= io_adcValues_77; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_78 <= io_adcValues_78; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_79 <= io_adcValues_79; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_80 <= io_adcValues_80; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_81 <= io_adcValues_81; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_82 <= io_adcValues_82; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_83 <= io_adcValues_83; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_84 <= io_adcValues_84; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_85 <= io_adcValues_85; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_86 <= io_adcValues_86; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_87 <= io_adcValues_87; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_88 <= io_adcValues_88; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_89 <= io_adcValues_89; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_90 <= io_adcValues_90; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_91 <= io_adcValues_91; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_92 <= io_adcValues_92; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_93 <= io_adcValues_93; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_94 <= io_adcValues_94; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_95 <= io_adcValues_95; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_96 <= io_adcValues_96; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_97 <= io_adcValues_97; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_98 <= io_adcValues_98; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_99 <= io_adcValues_99; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_100 <= io_adcValues_100; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_101 <= io_adcValues_101; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_102 <= io_adcValues_102; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_103 <= io_adcValues_103; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_104 <= io_adcValues_104; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_105 <= io_adcValues_105; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_106 <= io_adcValues_106; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_107 <= io_adcValues_107; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_108 <= io_adcValues_108; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_109 <= io_adcValues_109; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_110 <= io_adcValues_110; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_111 <= io_adcValues_111; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_112 <= io_adcValues_112; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_113 <= io_adcValues_113; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_114 <= io_adcValues_114; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_115 <= io_adcValues_115; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_116 <= io_adcValues_116; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_117 <= io_adcValues_117; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_118 <= io_adcValues_118; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_119 <= io_adcValues_119; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_120 <= io_adcValues_120; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_121 <= io_adcValues_121; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_122 <= io_adcValues_122; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_123 <= io_adcValues_123; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_124 <= io_adcValues_124; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_125 <= io_adcValues_125; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_126 <= io_adcValues_126; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hd == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_13_127 <= io_adcValues_127; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_0 <= io_adcValues_0; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_1 <= io_adcValues_1; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_2 <= io_adcValues_2; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_3 <= io_adcValues_3; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_4 <= io_adcValues_4; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_5 <= io_adcValues_5; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_6 <= io_adcValues_6; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_7 <= io_adcValues_7; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_8 <= io_adcValues_8; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_9 <= io_adcValues_9; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_10 <= io_adcValues_10; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_11 <= io_adcValues_11; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_12 <= io_adcValues_12; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_13 <= io_adcValues_13; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_14 <= io_adcValues_14; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_15 <= io_adcValues_15; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_16 <= io_adcValues_16; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_17 <= io_adcValues_17; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_18 <= io_adcValues_18; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_19 <= io_adcValues_19; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_20 <= io_adcValues_20; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_21 <= io_adcValues_21; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_22 <= io_adcValues_22; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_23 <= io_adcValues_23; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_24 <= io_adcValues_24; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_25 <= io_adcValues_25; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_26 <= io_adcValues_26; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_27 <= io_adcValues_27; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_28 <= io_adcValues_28; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_29 <= io_adcValues_29; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_30 <= io_adcValues_30; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_31 <= io_adcValues_31; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_32 <= io_adcValues_32; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_33 <= io_adcValues_33; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_34 <= io_adcValues_34; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_35 <= io_adcValues_35; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_36 <= io_adcValues_36; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_37 <= io_adcValues_37; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_38 <= io_adcValues_38; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_39 <= io_adcValues_39; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_40 <= io_adcValues_40; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_41 <= io_adcValues_41; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_42 <= io_adcValues_42; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_43 <= io_adcValues_43; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_44 <= io_adcValues_44; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_45 <= io_adcValues_45; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_46 <= io_adcValues_46; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_47 <= io_adcValues_47; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_48 <= io_adcValues_48; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_49 <= io_adcValues_49; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_50 <= io_adcValues_50; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_51 <= io_adcValues_51; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_52 <= io_adcValues_52; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_53 <= io_adcValues_53; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_54 <= io_adcValues_54; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_55 <= io_adcValues_55; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_56 <= io_adcValues_56; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_57 <= io_adcValues_57; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_58 <= io_adcValues_58; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_59 <= io_adcValues_59; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_60 <= io_adcValues_60; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_61 <= io_adcValues_61; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_62 <= io_adcValues_62; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_63 <= io_adcValues_63; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_64 <= io_adcValues_64; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_65 <= io_adcValues_65; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_66 <= io_adcValues_66; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_67 <= io_adcValues_67; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_68 <= io_adcValues_68; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_69 <= io_adcValues_69; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_70 <= io_adcValues_70; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_71 <= io_adcValues_71; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_72 <= io_adcValues_72; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_73 <= io_adcValues_73; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_74 <= io_adcValues_74; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_75 <= io_adcValues_75; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_76 <= io_adcValues_76; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_77 <= io_adcValues_77; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_78 <= io_adcValues_78; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_79 <= io_adcValues_79; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_80 <= io_adcValues_80; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_81 <= io_adcValues_81; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_82 <= io_adcValues_82; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_83 <= io_adcValues_83; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_84 <= io_adcValues_84; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_85 <= io_adcValues_85; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_86 <= io_adcValues_86; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_87 <= io_adcValues_87; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_88 <= io_adcValues_88; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_89 <= io_adcValues_89; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_90 <= io_adcValues_90; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_91 <= io_adcValues_91; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_92 <= io_adcValues_92; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_93 <= io_adcValues_93; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_94 <= io_adcValues_94; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_95 <= io_adcValues_95; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_96 <= io_adcValues_96; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_97 <= io_adcValues_97; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_98 <= io_adcValues_98; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_99 <= io_adcValues_99; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_100 <= io_adcValues_100; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_101 <= io_adcValues_101; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_102 <= io_adcValues_102; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_103 <= io_adcValues_103; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_104 <= io_adcValues_104; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_105 <= io_adcValues_105; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_106 <= io_adcValues_106; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_107 <= io_adcValues_107; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_108 <= io_adcValues_108; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_109 <= io_adcValues_109; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_110 <= io_adcValues_110; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_111 <= io_adcValues_111; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_112 <= io_adcValues_112; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_113 <= io_adcValues_113; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_114 <= io_adcValues_114; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_115 <= io_adcValues_115; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_116 <= io_adcValues_116; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_117 <= io_adcValues_117; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_118 <= io_adcValues_118; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_119 <= io_adcValues_119; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_120 <= io_adcValues_120; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_121 <= io_adcValues_121; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_122 <= io_adcValues_122; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_123 <= io_adcValues_123; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_124 <= io_adcValues_124; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_125 <= io_adcValues_125; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_126 <= io_adcValues_126; // @[BufferAMSNew.scala 24:28]
    end
    if (4'he == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_14_127 <= io_adcValues_127; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_0 <= io_adcValues_0; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_1 <= io_adcValues_1; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_2 <= io_adcValues_2; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_3 <= io_adcValues_3; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_4 <= io_adcValues_4; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_5 <= io_adcValues_5; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_6 <= io_adcValues_6; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_7 <= io_adcValues_7; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_8 <= io_adcValues_8; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_9 <= io_adcValues_9; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_10 <= io_adcValues_10; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_11 <= io_adcValues_11; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_12 <= io_adcValues_12; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_13 <= io_adcValues_13; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_14 <= io_adcValues_14; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_15 <= io_adcValues_15; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_16 <= io_adcValues_16; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_17 <= io_adcValues_17; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_18 <= io_adcValues_18; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_19 <= io_adcValues_19; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_20 <= io_adcValues_20; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_21 <= io_adcValues_21; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_22 <= io_adcValues_22; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_23 <= io_adcValues_23; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_24 <= io_adcValues_24; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_25 <= io_adcValues_25; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_26 <= io_adcValues_26; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_27 <= io_adcValues_27; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_28 <= io_adcValues_28; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_29 <= io_adcValues_29; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_30 <= io_adcValues_30; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_31 <= io_adcValues_31; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_32 <= io_adcValues_32; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_33 <= io_adcValues_33; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_34 <= io_adcValues_34; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_35 <= io_adcValues_35; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_36 <= io_adcValues_36; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_37 <= io_adcValues_37; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_38 <= io_adcValues_38; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_39 <= io_adcValues_39; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_40 <= io_adcValues_40; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_41 <= io_adcValues_41; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_42 <= io_adcValues_42; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_43 <= io_adcValues_43; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_44 <= io_adcValues_44; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_45 <= io_adcValues_45; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_46 <= io_adcValues_46; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_47 <= io_adcValues_47; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_48 <= io_adcValues_48; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_49 <= io_adcValues_49; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_50 <= io_adcValues_50; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_51 <= io_adcValues_51; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_52 <= io_adcValues_52; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_53 <= io_adcValues_53; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_54 <= io_adcValues_54; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_55 <= io_adcValues_55; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_56 <= io_adcValues_56; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_57 <= io_adcValues_57; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_58 <= io_adcValues_58; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_59 <= io_adcValues_59; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_60 <= io_adcValues_60; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_61 <= io_adcValues_61; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_62 <= io_adcValues_62; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_63 <= io_adcValues_63; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_64 <= io_adcValues_64; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_65 <= io_adcValues_65; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_66 <= io_adcValues_66; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_67 <= io_adcValues_67; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_68 <= io_adcValues_68; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_69 <= io_adcValues_69; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_70 <= io_adcValues_70; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_71 <= io_adcValues_71; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_72 <= io_adcValues_72; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_73 <= io_adcValues_73; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_74 <= io_adcValues_74; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_75 <= io_adcValues_75; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_76 <= io_adcValues_76; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_77 <= io_adcValues_77; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_78 <= io_adcValues_78; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_79 <= io_adcValues_79; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_80 <= io_adcValues_80; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_81 <= io_adcValues_81; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_82 <= io_adcValues_82; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_83 <= io_adcValues_83; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_84 <= io_adcValues_84; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_85 <= io_adcValues_85; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_86 <= io_adcValues_86; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_87 <= io_adcValues_87; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_88 <= io_adcValues_88; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_89 <= io_adcValues_89; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_90 <= io_adcValues_90; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_91 <= io_adcValues_91; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_92 <= io_adcValues_92; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_93 <= io_adcValues_93; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_94 <= io_adcValues_94; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_95 <= io_adcValues_95; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_96 <= io_adcValues_96; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_97 <= io_adcValues_97; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_98 <= io_adcValues_98; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_99 <= io_adcValues_99; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_100 <= io_adcValues_100; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_101 <= io_adcValues_101; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_102 <= io_adcValues_102; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_103 <= io_adcValues_103; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_104 <= io_adcValues_104; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_105 <= io_adcValues_105; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_106 <= io_adcValues_106; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_107 <= io_adcValues_107; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_108 <= io_adcValues_108; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_109 <= io_adcValues_109; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_110 <= io_adcValues_110; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_111 <= io_adcValues_111; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_112 <= io_adcValues_112; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_113 <= io_adcValues_113; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_114 <= io_adcValues_114; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_115 <= io_adcValues_115; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_116 <= io_adcValues_116; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_117 <= io_adcValues_117; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_118 <= io_adcValues_118; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_119 <= io_adcValues_119; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_120 <= io_adcValues_120; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_121 <= io_adcValues_121; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_122 <= io_adcValues_122; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_123 <= io_adcValues_123; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_124 <= io_adcValues_124; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_125 <= io_adcValues_125; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_126 <= io_adcValues_126; // @[BufferAMSNew.scala 24:28]
    end
    if (4'hf == lineCounter) begin // @[BufferAMSNew.scala 24:28]
      frameBuffer_15_127 <= io_adcValues_127; // @[BufferAMSNew.scala 24:28]
    end
    if (reset) begin // @[BufferAMSNew.scala 21:28]
      lineCounter <= 4'h0; // @[BufferAMSNew.scala 21:28]
    end else if (lineCounter == 4'hf) begin // @[BufferAMSNew.scala 28:30]
      lineCounter <= 4'h0; // @[BufferAMSNew.scala 29:17]
    end else begin
      lineCounter <= _lineCounter_T_1; // @[BufferAMSNew.scala 33:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  zeroAccumulators_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  zeroAccumulators_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  zeroAccumulators_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  zeroAccumulators_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  zeroAccumulators_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  zeroAccumulators_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  zeroAccumulators_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  zeroAccumulators_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  indexAccumulators_0 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  indexAccumulators_1 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  indexAccumulators_2 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  indexAccumulators_3 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  indexAccumulators_4 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  indexAccumulators_5 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  indexAccumulators_6 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  indexAccumulators_7 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  frameBuffer_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  frameBuffer_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  frameBuffer_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  frameBuffer_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  frameBuffer_0_4 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  frameBuffer_0_5 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  frameBuffer_0_6 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  frameBuffer_0_7 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  frameBuffer_0_8 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  frameBuffer_0_9 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  frameBuffer_0_10 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  frameBuffer_0_11 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  frameBuffer_0_12 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  frameBuffer_0_13 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  frameBuffer_0_14 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  frameBuffer_0_15 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  frameBuffer_0_16 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  frameBuffer_0_17 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  frameBuffer_0_18 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  frameBuffer_0_19 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  frameBuffer_0_20 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  frameBuffer_0_21 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  frameBuffer_0_22 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  frameBuffer_0_23 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  frameBuffer_0_24 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  frameBuffer_0_25 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  frameBuffer_0_26 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  frameBuffer_0_27 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  frameBuffer_0_28 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  frameBuffer_0_29 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  frameBuffer_0_30 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  frameBuffer_0_31 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  frameBuffer_0_32 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  frameBuffer_0_33 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  frameBuffer_0_34 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  frameBuffer_0_35 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  frameBuffer_0_36 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  frameBuffer_0_37 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  frameBuffer_0_38 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  frameBuffer_0_39 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  frameBuffer_0_40 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  frameBuffer_0_41 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  frameBuffer_0_42 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  frameBuffer_0_43 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  frameBuffer_0_44 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  frameBuffer_0_45 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  frameBuffer_0_46 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  frameBuffer_0_47 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  frameBuffer_0_48 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  frameBuffer_0_49 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  frameBuffer_0_50 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  frameBuffer_0_51 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  frameBuffer_0_52 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  frameBuffer_0_53 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  frameBuffer_0_54 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  frameBuffer_0_55 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  frameBuffer_0_56 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  frameBuffer_0_57 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  frameBuffer_0_58 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  frameBuffer_0_59 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  frameBuffer_0_60 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  frameBuffer_0_61 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  frameBuffer_0_62 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  frameBuffer_0_63 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  frameBuffer_0_64 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  frameBuffer_0_65 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  frameBuffer_0_66 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  frameBuffer_0_67 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  frameBuffer_0_68 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  frameBuffer_0_69 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  frameBuffer_0_70 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  frameBuffer_0_71 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  frameBuffer_0_72 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  frameBuffer_0_73 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  frameBuffer_0_74 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  frameBuffer_0_75 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  frameBuffer_0_76 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  frameBuffer_0_77 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  frameBuffer_0_78 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  frameBuffer_0_79 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  frameBuffer_0_80 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  frameBuffer_0_81 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  frameBuffer_0_82 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  frameBuffer_0_83 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  frameBuffer_0_84 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  frameBuffer_0_85 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  frameBuffer_0_86 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  frameBuffer_0_87 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  frameBuffer_0_88 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  frameBuffer_0_89 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  frameBuffer_0_90 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  frameBuffer_0_91 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  frameBuffer_0_92 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  frameBuffer_0_93 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  frameBuffer_0_94 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  frameBuffer_0_95 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  frameBuffer_0_96 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  frameBuffer_0_97 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  frameBuffer_0_98 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  frameBuffer_0_99 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  frameBuffer_0_100 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  frameBuffer_0_101 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  frameBuffer_0_102 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  frameBuffer_0_103 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  frameBuffer_0_104 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  frameBuffer_0_105 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  frameBuffer_0_106 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  frameBuffer_0_107 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  frameBuffer_0_108 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  frameBuffer_0_109 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  frameBuffer_0_110 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  frameBuffer_0_111 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  frameBuffer_0_112 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  frameBuffer_0_113 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  frameBuffer_0_114 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  frameBuffer_0_115 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  frameBuffer_0_116 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  frameBuffer_0_117 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  frameBuffer_0_118 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  frameBuffer_0_119 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  frameBuffer_0_120 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  frameBuffer_0_121 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  frameBuffer_0_122 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  frameBuffer_0_123 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  frameBuffer_0_124 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  frameBuffer_0_125 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  frameBuffer_0_126 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  frameBuffer_0_127 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  frameBuffer_1_0 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  frameBuffer_1_1 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  frameBuffer_1_2 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  frameBuffer_1_3 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  frameBuffer_1_4 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  frameBuffer_1_5 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  frameBuffer_1_6 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  frameBuffer_1_7 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  frameBuffer_1_8 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  frameBuffer_1_9 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  frameBuffer_1_10 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  frameBuffer_1_11 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  frameBuffer_1_12 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  frameBuffer_1_13 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  frameBuffer_1_14 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  frameBuffer_1_15 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  frameBuffer_1_16 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  frameBuffer_1_17 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  frameBuffer_1_18 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  frameBuffer_1_19 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  frameBuffer_1_20 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  frameBuffer_1_21 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  frameBuffer_1_22 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  frameBuffer_1_23 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  frameBuffer_1_24 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  frameBuffer_1_25 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  frameBuffer_1_26 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  frameBuffer_1_27 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  frameBuffer_1_28 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  frameBuffer_1_29 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  frameBuffer_1_30 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  frameBuffer_1_31 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  frameBuffer_1_32 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  frameBuffer_1_33 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  frameBuffer_1_34 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  frameBuffer_1_35 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  frameBuffer_1_36 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  frameBuffer_1_37 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  frameBuffer_1_38 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  frameBuffer_1_39 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  frameBuffer_1_40 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  frameBuffer_1_41 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  frameBuffer_1_42 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  frameBuffer_1_43 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  frameBuffer_1_44 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  frameBuffer_1_45 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  frameBuffer_1_46 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  frameBuffer_1_47 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  frameBuffer_1_48 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  frameBuffer_1_49 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  frameBuffer_1_50 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  frameBuffer_1_51 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  frameBuffer_1_52 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  frameBuffer_1_53 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  frameBuffer_1_54 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  frameBuffer_1_55 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  frameBuffer_1_56 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  frameBuffer_1_57 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  frameBuffer_1_58 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  frameBuffer_1_59 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  frameBuffer_1_60 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  frameBuffer_1_61 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  frameBuffer_1_62 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  frameBuffer_1_63 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  frameBuffer_1_64 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  frameBuffer_1_65 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  frameBuffer_1_66 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  frameBuffer_1_67 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  frameBuffer_1_68 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  frameBuffer_1_69 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  frameBuffer_1_70 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  frameBuffer_1_71 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  frameBuffer_1_72 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  frameBuffer_1_73 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  frameBuffer_1_74 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  frameBuffer_1_75 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  frameBuffer_1_76 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  frameBuffer_1_77 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  frameBuffer_1_78 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  frameBuffer_1_79 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  frameBuffer_1_80 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  frameBuffer_1_81 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  frameBuffer_1_82 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  frameBuffer_1_83 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  frameBuffer_1_84 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  frameBuffer_1_85 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  frameBuffer_1_86 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  frameBuffer_1_87 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  frameBuffer_1_88 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  frameBuffer_1_89 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  frameBuffer_1_90 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  frameBuffer_1_91 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  frameBuffer_1_92 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  frameBuffer_1_93 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  frameBuffer_1_94 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  frameBuffer_1_95 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  frameBuffer_1_96 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  frameBuffer_1_97 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  frameBuffer_1_98 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  frameBuffer_1_99 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  frameBuffer_1_100 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  frameBuffer_1_101 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  frameBuffer_1_102 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  frameBuffer_1_103 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  frameBuffer_1_104 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  frameBuffer_1_105 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  frameBuffer_1_106 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  frameBuffer_1_107 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  frameBuffer_1_108 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  frameBuffer_1_109 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  frameBuffer_1_110 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  frameBuffer_1_111 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  frameBuffer_1_112 = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  frameBuffer_1_113 = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  frameBuffer_1_114 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  frameBuffer_1_115 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  frameBuffer_1_116 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  frameBuffer_1_117 = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  frameBuffer_1_118 = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  frameBuffer_1_119 = _RAND_263[7:0];
  _RAND_264 = {1{`RANDOM}};
  frameBuffer_1_120 = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  frameBuffer_1_121 = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  frameBuffer_1_122 = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  frameBuffer_1_123 = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  frameBuffer_1_124 = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  frameBuffer_1_125 = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  frameBuffer_1_126 = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  frameBuffer_1_127 = _RAND_271[7:0];
  _RAND_272 = {1{`RANDOM}};
  frameBuffer_2_0 = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  frameBuffer_2_1 = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  frameBuffer_2_2 = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  frameBuffer_2_3 = _RAND_275[7:0];
  _RAND_276 = {1{`RANDOM}};
  frameBuffer_2_4 = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  frameBuffer_2_5 = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  frameBuffer_2_6 = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  frameBuffer_2_7 = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  frameBuffer_2_8 = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  frameBuffer_2_9 = _RAND_281[7:0];
  _RAND_282 = {1{`RANDOM}};
  frameBuffer_2_10 = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  frameBuffer_2_11 = _RAND_283[7:0];
  _RAND_284 = {1{`RANDOM}};
  frameBuffer_2_12 = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  frameBuffer_2_13 = _RAND_285[7:0];
  _RAND_286 = {1{`RANDOM}};
  frameBuffer_2_14 = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  frameBuffer_2_15 = _RAND_287[7:0];
  _RAND_288 = {1{`RANDOM}};
  frameBuffer_2_16 = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  frameBuffer_2_17 = _RAND_289[7:0];
  _RAND_290 = {1{`RANDOM}};
  frameBuffer_2_18 = _RAND_290[7:0];
  _RAND_291 = {1{`RANDOM}};
  frameBuffer_2_19 = _RAND_291[7:0];
  _RAND_292 = {1{`RANDOM}};
  frameBuffer_2_20 = _RAND_292[7:0];
  _RAND_293 = {1{`RANDOM}};
  frameBuffer_2_21 = _RAND_293[7:0];
  _RAND_294 = {1{`RANDOM}};
  frameBuffer_2_22 = _RAND_294[7:0];
  _RAND_295 = {1{`RANDOM}};
  frameBuffer_2_23 = _RAND_295[7:0];
  _RAND_296 = {1{`RANDOM}};
  frameBuffer_2_24 = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  frameBuffer_2_25 = _RAND_297[7:0];
  _RAND_298 = {1{`RANDOM}};
  frameBuffer_2_26 = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  frameBuffer_2_27 = _RAND_299[7:0];
  _RAND_300 = {1{`RANDOM}};
  frameBuffer_2_28 = _RAND_300[7:0];
  _RAND_301 = {1{`RANDOM}};
  frameBuffer_2_29 = _RAND_301[7:0];
  _RAND_302 = {1{`RANDOM}};
  frameBuffer_2_30 = _RAND_302[7:0];
  _RAND_303 = {1{`RANDOM}};
  frameBuffer_2_31 = _RAND_303[7:0];
  _RAND_304 = {1{`RANDOM}};
  frameBuffer_2_32 = _RAND_304[7:0];
  _RAND_305 = {1{`RANDOM}};
  frameBuffer_2_33 = _RAND_305[7:0];
  _RAND_306 = {1{`RANDOM}};
  frameBuffer_2_34 = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  frameBuffer_2_35 = _RAND_307[7:0];
  _RAND_308 = {1{`RANDOM}};
  frameBuffer_2_36 = _RAND_308[7:0];
  _RAND_309 = {1{`RANDOM}};
  frameBuffer_2_37 = _RAND_309[7:0];
  _RAND_310 = {1{`RANDOM}};
  frameBuffer_2_38 = _RAND_310[7:0];
  _RAND_311 = {1{`RANDOM}};
  frameBuffer_2_39 = _RAND_311[7:0];
  _RAND_312 = {1{`RANDOM}};
  frameBuffer_2_40 = _RAND_312[7:0];
  _RAND_313 = {1{`RANDOM}};
  frameBuffer_2_41 = _RAND_313[7:0];
  _RAND_314 = {1{`RANDOM}};
  frameBuffer_2_42 = _RAND_314[7:0];
  _RAND_315 = {1{`RANDOM}};
  frameBuffer_2_43 = _RAND_315[7:0];
  _RAND_316 = {1{`RANDOM}};
  frameBuffer_2_44 = _RAND_316[7:0];
  _RAND_317 = {1{`RANDOM}};
  frameBuffer_2_45 = _RAND_317[7:0];
  _RAND_318 = {1{`RANDOM}};
  frameBuffer_2_46 = _RAND_318[7:0];
  _RAND_319 = {1{`RANDOM}};
  frameBuffer_2_47 = _RAND_319[7:0];
  _RAND_320 = {1{`RANDOM}};
  frameBuffer_2_48 = _RAND_320[7:0];
  _RAND_321 = {1{`RANDOM}};
  frameBuffer_2_49 = _RAND_321[7:0];
  _RAND_322 = {1{`RANDOM}};
  frameBuffer_2_50 = _RAND_322[7:0];
  _RAND_323 = {1{`RANDOM}};
  frameBuffer_2_51 = _RAND_323[7:0];
  _RAND_324 = {1{`RANDOM}};
  frameBuffer_2_52 = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  frameBuffer_2_53 = _RAND_325[7:0];
  _RAND_326 = {1{`RANDOM}};
  frameBuffer_2_54 = _RAND_326[7:0];
  _RAND_327 = {1{`RANDOM}};
  frameBuffer_2_55 = _RAND_327[7:0];
  _RAND_328 = {1{`RANDOM}};
  frameBuffer_2_56 = _RAND_328[7:0];
  _RAND_329 = {1{`RANDOM}};
  frameBuffer_2_57 = _RAND_329[7:0];
  _RAND_330 = {1{`RANDOM}};
  frameBuffer_2_58 = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  frameBuffer_2_59 = _RAND_331[7:0];
  _RAND_332 = {1{`RANDOM}};
  frameBuffer_2_60 = _RAND_332[7:0];
  _RAND_333 = {1{`RANDOM}};
  frameBuffer_2_61 = _RAND_333[7:0];
  _RAND_334 = {1{`RANDOM}};
  frameBuffer_2_62 = _RAND_334[7:0];
  _RAND_335 = {1{`RANDOM}};
  frameBuffer_2_63 = _RAND_335[7:0];
  _RAND_336 = {1{`RANDOM}};
  frameBuffer_2_64 = _RAND_336[7:0];
  _RAND_337 = {1{`RANDOM}};
  frameBuffer_2_65 = _RAND_337[7:0];
  _RAND_338 = {1{`RANDOM}};
  frameBuffer_2_66 = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  frameBuffer_2_67 = _RAND_339[7:0];
  _RAND_340 = {1{`RANDOM}};
  frameBuffer_2_68 = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  frameBuffer_2_69 = _RAND_341[7:0];
  _RAND_342 = {1{`RANDOM}};
  frameBuffer_2_70 = _RAND_342[7:0];
  _RAND_343 = {1{`RANDOM}};
  frameBuffer_2_71 = _RAND_343[7:0];
  _RAND_344 = {1{`RANDOM}};
  frameBuffer_2_72 = _RAND_344[7:0];
  _RAND_345 = {1{`RANDOM}};
  frameBuffer_2_73 = _RAND_345[7:0];
  _RAND_346 = {1{`RANDOM}};
  frameBuffer_2_74 = _RAND_346[7:0];
  _RAND_347 = {1{`RANDOM}};
  frameBuffer_2_75 = _RAND_347[7:0];
  _RAND_348 = {1{`RANDOM}};
  frameBuffer_2_76 = _RAND_348[7:0];
  _RAND_349 = {1{`RANDOM}};
  frameBuffer_2_77 = _RAND_349[7:0];
  _RAND_350 = {1{`RANDOM}};
  frameBuffer_2_78 = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  frameBuffer_2_79 = _RAND_351[7:0];
  _RAND_352 = {1{`RANDOM}};
  frameBuffer_2_80 = _RAND_352[7:0];
  _RAND_353 = {1{`RANDOM}};
  frameBuffer_2_81 = _RAND_353[7:0];
  _RAND_354 = {1{`RANDOM}};
  frameBuffer_2_82 = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  frameBuffer_2_83 = _RAND_355[7:0];
  _RAND_356 = {1{`RANDOM}};
  frameBuffer_2_84 = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  frameBuffer_2_85 = _RAND_357[7:0];
  _RAND_358 = {1{`RANDOM}};
  frameBuffer_2_86 = _RAND_358[7:0];
  _RAND_359 = {1{`RANDOM}};
  frameBuffer_2_87 = _RAND_359[7:0];
  _RAND_360 = {1{`RANDOM}};
  frameBuffer_2_88 = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  frameBuffer_2_89 = _RAND_361[7:0];
  _RAND_362 = {1{`RANDOM}};
  frameBuffer_2_90 = _RAND_362[7:0];
  _RAND_363 = {1{`RANDOM}};
  frameBuffer_2_91 = _RAND_363[7:0];
  _RAND_364 = {1{`RANDOM}};
  frameBuffer_2_92 = _RAND_364[7:0];
  _RAND_365 = {1{`RANDOM}};
  frameBuffer_2_93 = _RAND_365[7:0];
  _RAND_366 = {1{`RANDOM}};
  frameBuffer_2_94 = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  frameBuffer_2_95 = _RAND_367[7:0];
  _RAND_368 = {1{`RANDOM}};
  frameBuffer_2_96 = _RAND_368[7:0];
  _RAND_369 = {1{`RANDOM}};
  frameBuffer_2_97 = _RAND_369[7:0];
  _RAND_370 = {1{`RANDOM}};
  frameBuffer_2_98 = _RAND_370[7:0];
  _RAND_371 = {1{`RANDOM}};
  frameBuffer_2_99 = _RAND_371[7:0];
  _RAND_372 = {1{`RANDOM}};
  frameBuffer_2_100 = _RAND_372[7:0];
  _RAND_373 = {1{`RANDOM}};
  frameBuffer_2_101 = _RAND_373[7:0];
  _RAND_374 = {1{`RANDOM}};
  frameBuffer_2_102 = _RAND_374[7:0];
  _RAND_375 = {1{`RANDOM}};
  frameBuffer_2_103 = _RAND_375[7:0];
  _RAND_376 = {1{`RANDOM}};
  frameBuffer_2_104 = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  frameBuffer_2_105 = _RAND_377[7:0];
  _RAND_378 = {1{`RANDOM}};
  frameBuffer_2_106 = _RAND_378[7:0];
  _RAND_379 = {1{`RANDOM}};
  frameBuffer_2_107 = _RAND_379[7:0];
  _RAND_380 = {1{`RANDOM}};
  frameBuffer_2_108 = _RAND_380[7:0];
  _RAND_381 = {1{`RANDOM}};
  frameBuffer_2_109 = _RAND_381[7:0];
  _RAND_382 = {1{`RANDOM}};
  frameBuffer_2_110 = _RAND_382[7:0];
  _RAND_383 = {1{`RANDOM}};
  frameBuffer_2_111 = _RAND_383[7:0];
  _RAND_384 = {1{`RANDOM}};
  frameBuffer_2_112 = _RAND_384[7:0];
  _RAND_385 = {1{`RANDOM}};
  frameBuffer_2_113 = _RAND_385[7:0];
  _RAND_386 = {1{`RANDOM}};
  frameBuffer_2_114 = _RAND_386[7:0];
  _RAND_387 = {1{`RANDOM}};
  frameBuffer_2_115 = _RAND_387[7:0];
  _RAND_388 = {1{`RANDOM}};
  frameBuffer_2_116 = _RAND_388[7:0];
  _RAND_389 = {1{`RANDOM}};
  frameBuffer_2_117 = _RAND_389[7:0];
  _RAND_390 = {1{`RANDOM}};
  frameBuffer_2_118 = _RAND_390[7:0];
  _RAND_391 = {1{`RANDOM}};
  frameBuffer_2_119 = _RAND_391[7:0];
  _RAND_392 = {1{`RANDOM}};
  frameBuffer_2_120 = _RAND_392[7:0];
  _RAND_393 = {1{`RANDOM}};
  frameBuffer_2_121 = _RAND_393[7:0];
  _RAND_394 = {1{`RANDOM}};
  frameBuffer_2_122 = _RAND_394[7:0];
  _RAND_395 = {1{`RANDOM}};
  frameBuffer_2_123 = _RAND_395[7:0];
  _RAND_396 = {1{`RANDOM}};
  frameBuffer_2_124 = _RAND_396[7:0];
  _RAND_397 = {1{`RANDOM}};
  frameBuffer_2_125 = _RAND_397[7:0];
  _RAND_398 = {1{`RANDOM}};
  frameBuffer_2_126 = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  frameBuffer_2_127 = _RAND_399[7:0];
  _RAND_400 = {1{`RANDOM}};
  frameBuffer_3_0 = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  frameBuffer_3_1 = _RAND_401[7:0];
  _RAND_402 = {1{`RANDOM}};
  frameBuffer_3_2 = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  frameBuffer_3_3 = _RAND_403[7:0];
  _RAND_404 = {1{`RANDOM}};
  frameBuffer_3_4 = _RAND_404[7:0];
  _RAND_405 = {1{`RANDOM}};
  frameBuffer_3_5 = _RAND_405[7:0];
  _RAND_406 = {1{`RANDOM}};
  frameBuffer_3_6 = _RAND_406[7:0];
  _RAND_407 = {1{`RANDOM}};
  frameBuffer_3_7 = _RAND_407[7:0];
  _RAND_408 = {1{`RANDOM}};
  frameBuffer_3_8 = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  frameBuffer_3_9 = _RAND_409[7:0];
  _RAND_410 = {1{`RANDOM}};
  frameBuffer_3_10 = _RAND_410[7:0];
  _RAND_411 = {1{`RANDOM}};
  frameBuffer_3_11 = _RAND_411[7:0];
  _RAND_412 = {1{`RANDOM}};
  frameBuffer_3_12 = _RAND_412[7:0];
  _RAND_413 = {1{`RANDOM}};
  frameBuffer_3_13 = _RAND_413[7:0];
  _RAND_414 = {1{`RANDOM}};
  frameBuffer_3_14 = _RAND_414[7:0];
  _RAND_415 = {1{`RANDOM}};
  frameBuffer_3_15 = _RAND_415[7:0];
  _RAND_416 = {1{`RANDOM}};
  frameBuffer_3_16 = _RAND_416[7:0];
  _RAND_417 = {1{`RANDOM}};
  frameBuffer_3_17 = _RAND_417[7:0];
  _RAND_418 = {1{`RANDOM}};
  frameBuffer_3_18 = _RAND_418[7:0];
  _RAND_419 = {1{`RANDOM}};
  frameBuffer_3_19 = _RAND_419[7:0];
  _RAND_420 = {1{`RANDOM}};
  frameBuffer_3_20 = _RAND_420[7:0];
  _RAND_421 = {1{`RANDOM}};
  frameBuffer_3_21 = _RAND_421[7:0];
  _RAND_422 = {1{`RANDOM}};
  frameBuffer_3_22 = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  frameBuffer_3_23 = _RAND_423[7:0];
  _RAND_424 = {1{`RANDOM}};
  frameBuffer_3_24 = _RAND_424[7:0];
  _RAND_425 = {1{`RANDOM}};
  frameBuffer_3_25 = _RAND_425[7:0];
  _RAND_426 = {1{`RANDOM}};
  frameBuffer_3_26 = _RAND_426[7:0];
  _RAND_427 = {1{`RANDOM}};
  frameBuffer_3_27 = _RAND_427[7:0];
  _RAND_428 = {1{`RANDOM}};
  frameBuffer_3_28 = _RAND_428[7:0];
  _RAND_429 = {1{`RANDOM}};
  frameBuffer_3_29 = _RAND_429[7:0];
  _RAND_430 = {1{`RANDOM}};
  frameBuffer_3_30 = _RAND_430[7:0];
  _RAND_431 = {1{`RANDOM}};
  frameBuffer_3_31 = _RAND_431[7:0];
  _RAND_432 = {1{`RANDOM}};
  frameBuffer_3_32 = _RAND_432[7:0];
  _RAND_433 = {1{`RANDOM}};
  frameBuffer_3_33 = _RAND_433[7:0];
  _RAND_434 = {1{`RANDOM}};
  frameBuffer_3_34 = _RAND_434[7:0];
  _RAND_435 = {1{`RANDOM}};
  frameBuffer_3_35 = _RAND_435[7:0];
  _RAND_436 = {1{`RANDOM}};
  frameBuffer_3_36 = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  frameBuffer_3_37 = _RAND_437[7:0];
  _RAND_438 = {1{`RANDOM}};
  frameBuffer_3_38 = _RAND_438[7:0];
  _RAND_439 = {1{`RANDOM}};
  frameBuffer_3_39 = _RAND_439[7:0];
  _RAND_440 = {1{`RANDOM}};
  frameBuffer_3_40 = _RAND_440[7:0];
  _RAND_441 = {1{`RANDOM}};
  frameBuffer_3_41 = _RAND_441[7:0];
  _RAND_442 = {1{`RANDOM}};
  frameBuffer_3_42 = _RAND_442[7:0];
  _RAND_443 = {1{`RANDOM}};
  frameBuffer_3_43 = _RAND_443[7:0];
  _RAND_444 = {1{`RANDOM}};
  frameBuffer_3_44 = _RAND_444[7:0];
  _RAND_445 = {1{`RANDOM}};
  frameBuffer_3_45 = _RAND_445[7:0];
  _RAND_446 = {1{`RANDOM}};
  frameBuffer_3_46 = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  frameBuffer_3_47 = _RAND_447[7:0];
  _RAND_448 = {1{`RANDOM}};
  frameBuffer_3_48 = _RAND_448[7:0];
  _RAND_449 = {1{`RANDOM}};
  frameBuffer_3_49 = _RAND_449[7:0];
  _RAND_450 = {1{`RANDOM}};
  frameBuffer_3_50 = _RAND_450[7:0];
  _RAND_451 = {1{`RANDOM}};
  frameBuffer_3_51 = _RAND_451[7:0];
  _RAND_452 = {1{`RANDOM}};
  frameBuffer_3_52 = _RAND_452[7:0];
  _RAND_453 = {1{`RANDOM}};
  frameBuffer_3_53 = _RAND_453[7:0];
  _RAND_454 = {1{`RANDOM}};
  frameBuffer_3_54 = _RAND_454[7:0];
  _RAND_455 = {1{`RANDOM}};
  frameBuffer_3_55 = _RAND_455[7:0];
  _RAND_456 = {1{`RANDOM}};
  frameBuffer_3_56 = _RAND_456[7:0];
  _RAND_457 = {1{`RANDOM}};
  frameBuffer_3_57 = _RAND_457[7:0];
  _RAND_458 = {1{`RANDOM}};
  frameBuffer_3_58 = _RAND_458[7:0];
  _RAND_459 = {1{`RANDOM}};
  frameBuffer_3_59 = _RAND_459[7:0];
  _RAND_460 = {1{`RANDOM}};
  frameBuffer_3_60 = _RAND_460[7:0];
  _RAND_461 = {1{`RANDOM}};
  frameBuffer_3_61 = _RAND_461[7:0];
  _RAND_462 = {1{`RANDOM}};
  frameBuffer_3_62 = _RAND_462[7:0];
  _RAND_463 = {1{`RANDOM}};
  frameBuffer_3_63 = _RAND_463[7:0];
  _RAND_464 = {1{`RANDOM}};
  frameBuffer_3_64 = _RAND_464[7:0];
  _RAND_465 = {1{`RANDOM}};
  frameBuffer_3_65 = _RAND_465[7:0];
  _RAND_466 = {1{`RANDOM}};
  frameBuffer_3_66 = _RAND_466[7:0];
  _RAND_467 = {1{`RANDOM}};
  frameBuffer_3_67 = _RAND_467[7:0];
  _RAND_468 = {1{`RANDOM}};
  frameBuffer_3_68 = _RAND_468[7:0];
  _RAND_469 = {1{`RANDOM}};
  frameBuffer_3_69 = _RAND_469[7:0];
  _RAND_470 = {1{`RANDOM}};
  frameBuffer_3_70 = _RAND_470[7:0];
  _RAND_471 = {1{`RANDOM}};
  frameBuffer_3_71 = _RAND_471[7:0];
  _RAND_472 = {1{`RANDOM}};
  frameBuffer_3_72 = _RAND_472[7:0];
  _RAND_473 = {1{`RANDOM}};
  frameBuffer_3_73 = _RAND_473[7:0];
  _RAND_474 = {1{`RANDOM}};
  frameBuffer_3_74 = _RAND_474[7:0];
  _RAND_475 = {1{`RANDOM}};
  frameBuffer_3_75 = _RAND_475[7:0];
  _RAND_476 = {1{`RANDOM}};
  frameBuffer_3_76 = _RAND_476[7:0];
  _RAND_477 = {1{`RANDOM}};
  frameBuffer_3_77 = _RAND_477[7:0];
  _RAND_478 = {1{`RANDOM}};
  frameBuffer_3_78 = _RAND_478[7:0];
  _RAND_479 = {1{`RANDOM}};
  frameBuffer_3_79 = _RAND_479[7:0];
  _RAND_480 = {1{`RANDOM}};
  frameBuffer_3_80 = _RAND_480[7:0];
  _RAND_481 = {1{`RANDOM}};
  frameBuffer_3_81 = _RAND_481[7:0];
  _RAND_482 = {1{`RANDOM}};
  frameBuffer_3_82 = _RAND_482[7:0];
  _RAND_483 = {1{`RANDOM}};
  frameBuffer_3_83 = _RAND_483[7:0];
  _RAND_484 = {1{`RANDOM}};
  frameBuffer_3_84 = _RAND_484[7:0];
  _RAND_485 = {1{`RANDOM}};
  frameBuffer_3_85 = _RAND_485[7:0];
  _RAND_486 = {1{`RANDOM}};
  frameBuffer_3_86 = _RAND_486[7:0];
  _RAND_487 = {1{`RANDOM}};
  frameBuffer_3_87 = _RAND_487[7:0];
  _RAND_488 = {1{`RANDOM}};
  frameBuffer_3_88 = _RAND_488[7:0];
  _RAND_489 = {1{`RANDOM}};
  frameBuffer_3_89 = _RAND_489[7:0];
  _RAND_490 = {1{`RANDOM}};
  frameBuffer_3_90 = _RAND_490[7:0];
  _RAND_491 = {1{`RANDOM}};
  frameBuffer_3_91 = _RAND_491[7:0];
  _RAND_492 = {1{`RANDOM}};
  frameBuffer_3_92 = _RAND_492[7:0];
  _RAND_493 = {1{`RANDOM}};
  frameBuffer_3_93 = _RAND_493[7:0];
  _RAND_494 = {1{`RANDOM}};
  frameBuffer_3_94 = _RAND_494[7:0];
  _RAND_495 = {1{`RANDOM}};
  frameBuffer_3_95 = _RAND_495[7:0];
  _RAND_496 = {1{`RANDOM}};
  frameBuffer_3_96 = _RAND_496[7:0];
  _RAND_497 = {1{`RANDOM}};
  frameBuffer_3_97 = _RAND_497[7:0];
  _RAND_498 = {1{`RANDOM}};
  frameBuffer_3_98 = _RAND_498[7:0];
  _RAND_499 = {1{`RANDOM}};
  frameBuffer_3_99 = _RAND_499[7:0];
  _RAND_500 = {1{`RANDOM}};
  frameBuffer_3_100 = _RAND_500[7:0];
  _RAND_501 = {1{`RANDOM}};
  frameBuffer_3_101 = _RAND_501[7:0];
  _RAND_502 = {1{`RANDOM}};
  frameBuffer_3_102 = _RAND_502[7:0];
  _RAND_503 = {1{`RANDOM}};
  frameBuffer_3_103 = _RAND_503[7:0];
  _RAND_504 = {1{`RANDOM}};
  frameBuffer_3_104 = _RAND_504[7:0];
  _RAND_505 = {1{`RANDOM}};
  frameBuffer_3_105 = _RAND_505[7:0];
  _RAND_506 = {1{`RANDOM}};
  frameBuffer_3_106 = _RAND_506[7:0];
  _RAND_507 = {1{`RANDOM}};
  frameBuffer_3_107 = _RAND_507[7:0];
  _RAND_508 = {1{`RANDOM}};
  frameBuffer_3_108 = _RAND_508[7:0];
  _RAND_509 = {1{`RANDOM}};
  frameBuffer_3_109 = _RAND_509[7:0];
  _RAND_510 = {1{`RANDOM}};
  frameBuffer_3_110 = _RAND_510[7:0];
  _RAND_511 = {1{`RANDOM}};
  frameBuffer_3_111 = _RAND_511[7:0];
  _RAND_512 = {1{`RANDOM}};
  frameBuffer_3_112 = _RAND_512[7:0];
  _RAND_513 = {1{`RANDOM}};
  frameBuffer_3_113 = _RAND_513[7:0];
  _RAND_514 = {1{`RANDOM}};
  frameBuffer_3_114 = _RAND_514[7:0];
  _RAND_515 = {1{`RANDOM}};
  frameBuffer_3_115 = _RAND_515[7:0];
  _RAND_516 = {1{`RANDOM}};
  frameBuffer_3_116 = _RAND_516[7:0];
  _RAND_517 = {1{`RANDOM}};
  frameBuffer_3_117 = _RAND_517[7:0];
  _RAND_518 = {1{`RANDOM}};
  frameBuffer_3_118 = _RAND_518[7:0];
  _RAND_519 = {1{`RANDOM}};
  frameBuffer_3_119 = _RAND_519[7:0];
  _RAND_520 = {1{`RANDOM}};
  frameBuffer_3_120 = _RAND_520[7:0];
  _RAND_521 = {1{`RANDOM}};
  frameBuffer_3_121 = _RAND_521[7:0];
  _RAND_522 = {1{`RANDOM}};
  frameBuffer_3_122 = _RAND_522[7:0];
  _RAND_523 = {1{`RANDOM}};
  frameBuffer_3_123 = _RAND_523[7:0];
  _RAND_524 = {1{`RANDOM}};
  frameBuffer_3_124 = _RAND_524[7:0];
  _RAND_525 = {1{`RANDOM}};
  frameBuffer_3_125 = _RAND_525[7:0];
  _RAND_526 = {1{`RANDOM}};
  frameBuffer_3_126 = _RAND_526[7:0];
  _RAND_527 = {1{`RANDOM}};
  frameBuffer_3_127 = _RAND_527[7:0];
  _RAND_528 = {1{`RANDOM}};
  frameBuffer_4_0 = _RAND_528[7:0];
  _RAND_529 = {1{`RANDOM}};
  frameBuffer_4_1 = _RAND_529[7:0];
  _RAND_530 = {1{`RANDOM}};
  frameBuffer_4_2 = _RAND_530[7:0];
  _RAND_531 = {1{`RANDOM}};
  frameBuffer_4_3 = _RAND_531[7:0];
  _RAND_532 = {1{`RANDOM}};
  frameBuffer_4_4 = _RAND_532[7:0];
  _RAND_533 = {1{`RANDOM}};
  frameBuffer_4_5 = _RAND_533[7:0];
  _RAND_534 = {1{`RANDOM}};
  frameBuffer_4_6 = _RAND_534[7:0];
  _RAND_535 = {1{`RANDOM}};
  frameBuffer_4_7 = _RAND_535[7:0];
  _RAND_536 = {1{`RANDOM}};
  frameBuffer_4_8 = _RAND_536[7:0];
  _RAND_537 = {1{`RANDOM}};
  frameBuffer_4_9 = _RAND_537[7:0];
  _RAND_538 = {1{`RANDOM}};
  frameBuffer_4_10 = _RAND_538[7:0];
  _RAND_539 = {1{`RANDOM}};
  frameBuffer_4_11 = _RAND_539[7:0];
  _RAND_540 = {1{`RANDOM}};
  frameBuffer_4_12 = _RAND_540[7:0];
  _RAND_541 = {1{`RANDOM}};
  frameBuffer_4_13 = _RAND_541[7:0];
  _RAND_542 = {1{`RANDOM}};
  frameBuffer_4_14 = _RAND_542[7:0];
  _RAND_543 = {1{`RANDOM}};
  frameBuffer_4_15 = _RAND_543[7:0];
  _RAND_544 = {1{`RANDOM}};
  frameBuffer_4_16 = _RAND_544[7:0];
  _RAND_545 = {1{`RANDOM}};
  frameBuffer_4_17 = _RAND_545[7:0];
  _RAND_546 = {1{`RANDOM}};
  frameBuffer_4_18 = _RAND_546[7:0];
  _RAND_547 = {1{`RANDOM}};
  frameBuffer_4_19 = _RAND_547[7:0];
  _RAND_548 = {1{`RANDOM}};
  frameBuffer_4_20 = _RAND_548[7:0];
  _RAND_549 = {1{`RANDOM}};
  frameBuffer_4_21 = _RAND_549[7:0];
  _RAND_550 = {1{`RANDOM}};
  frameBuffer_4_22 = _RAND_550[7:0];
  _RAND_551 = {1{`RANDOM}};
  frameBuffer_4_23 = _RAND_551[7:0];
  _RAND_552 = {1{`RANDOM}};
  frameBuffer_4_24 = _RAND_552[7:0];
  _RAND_553 = {1{`RANDOM}};
  frameBuffer_4_25 = _RAND_553[7:0];
  _RAND_554 = {1{`RANDOM}};
  frameBuffer_4_26 = _RAND_554[7:0];
  _RAND_555 = {1{`RANDOM}};
  frameBuffer_4_27 = _RAND_555[7:0];
  _RAND_556 = {1{`RANDOM}};
  frameBuffer_4_28 = _RAND_556[7:0];
  _RAND_557 = {1{`RANDOM}};
  frameBuffer_4_29 = _RAND_557[7:0];
  _RAND_558 = {1{`RANDOM}};
  frameBuffer_4_30 = _RAND_558[7:0];
  _RAND_559 = {1{`RANDOM}};
  frameBuffer_4_31 = _RAND_559[7:0];
  _RAND_560 = {1{`RANDOM}};
  frameBuffer_4_32 = _RAND_560[7:0];
  _RAND_561 = {1{`RANDOM}};
  frameBuffer_4_33 = _RAND_561[7:0];
  _RAND_562 = {1{`RANDOM}};
  frameBuffer_4_34 = _RAND_562[7:0];
  _RAND_563 = {1{`RANDOM}};
  frameBuffer_4_35 = _RAND_563[7:0];
  _RAND_564 = {1{`RANDOM}};
  frameBuffer_4_36 = _RAND_564[7:0];
  _RAND_565 = {1{`RANDOM}};
  frameBuffer_4_37 = _RAND_565[7:0];
  _RAND_566 = {1{`RANDOM}};
  frameBuffer_4_38 = _RAND_566[7:0];
  _RAND_567 = {1{`RANDOM}};
  frameBuffer_4_39 = _RAND_567[7:0];
  _RAND_568 = {1{`RANDOM}};
  frameBuffer_4_40 = _RAND_568[7:0];
  _RAND_569 = {1{`RANDOM}};
  frameBuffer_4_41 = _RAND_569[7:0];
  _RAND_570 = {1{`RANDOM}};
  frameBuffer_4_42 = _RAND_570[7:0];
  _RAND_571 = {1{`RANDOM}};
  frameBuffer_4_43 = _RAND_571[7:0];
  _RAND_572 = {1{`RANDOM}};
  frameBuffer_4_44 = _RAND_572[7:0];
  _RAND_573 = {1{`RANDOM}};
  frameBuffer_4_45 = _RAND_573[7:0];
  _RAND_574 = {1{`RANDOM}};
  frameBuffer_4_46 = _RAND_574[7:0];
  _RAND_575 = {1{`RANDOM}};
  frameBuffer_4_47 = _RAND_575[7:0];
  _RAND_576 = {1{`RANDOM}};
  frameBuffer_4_48 = _RAND_576[7:0];
  _RAND_577 = {1{`RANDOM}};
  frameBuffer_4_49 = _RAND_577[7:0];
  _RAND_578 = {1{`RANDOM}};
  frameBuffer_4_50 = _RAND_578[7:0];
  _RAND_579 = {1{`RANDOM}};
  frameBuffer_4_51 = _RAND_579[7:0];
  _RAND_580 = {1{`RANDOM}};
  frameBuffer_4_52 = _RAND_580[7:0];
  _RAND_581 = {1{`RANDOM}};
  frameBuffer_4_53 = _RAND_581[7:0];
  _RAND_582 = {1{`RANDOM}};
  frameBuffer_4_54 = _RAND_582[7:0];
  _RAND_583 = {1{`RANDOM}};
  frameBuffer_4_55 = _RAND_583[7:0];
  _RAND_584 = {1{`RANDOM}};
  frameBuffer_4_56 = _RAND_584[7:0];
  _RAND_585 = {1{`RANDOM}};
  frameBuffer_4_57 = _RAND_585[7:0];
  _RAND_586 = {1{`RANDOM}};
  frameBuffer_4_58 = _RAND_586[7:0];
  _RAND_587 = {1{`RANDOM}};
  frameBuffer_4_59 = _RAND_587[7:0];
  _RAND_588 = {1{`RANDOM}};
  frameBuffer_4_60 = _RAND_588[7:0];
  _RAND_589 = {1{`RANDOM}};
  frameBuffer_4_61 = _RAND_589[7:0];
  _RAND_590 = {1{`RANDOM}};
  frameBuffer_4_62 = _RAND_590[7:0];
  _RAND_591 = {1{`RANDOM}};
  frameBuffer_4_63 = _RAND_591[7:0];
  _RAND_592 = {1{`RANDOM}};
  frameBuffer_4_64 = _RAND_592[7:0];
  _RAND_593 = {1{`RANDOM}};
  frameBuffer_4_65 = _RAND_593[7:0];
  _RAND_594 = {1{`RANDOM}};
  frameBuffer_4_66 = _RAND_594[7:0];
  _RAND_595 = {1{`RANDOM}};
  frameBuffer_4_67 = _RAND_595[7:0];
  _RAND_596 = {1{`RANDOM}};
  frameBuffer_4_68 = _RAND_596[7:0];
  _RAND_597 = {1{`RANDOM}};
  frameBuffer_4_69 = _RAND_597[7:0];
  _RAND_598 = {1{`RANDOM}};
  frameBuffer_4_70 = _RAND_598[7:0];
  _RAND_599 = {1{`RANDOM}};
  frameBuffer_4_71 = _RAND_599[7:0];
  _RAND_600 = {1{`RANDOM}};
  frameBuffer_4_72 = _RAND_600[7:0];
  _RAND_601 = {1{`RANDOM}};
  frameBuffer_4_73 = _RAND_601[7:0];
  _RAND_602 = {1{`RANDOM}};
  frameBuffer_4_74 = _RAND_602[7:0];
  _RAND_603 = {1{`RANDOM}};
  frameBuffer_4_75 = _RAND_603[7:0];
  _RAND_604 = {1{`RANDOM}};
  frameBuffer_4_76 = _RAND_604[7:0];
  _RAND_605 = {1{`RANDOM}};
  frameBuffer_4_77 = _RAND_605[7:0];
  _RAND_606 = {1{`RANDOM}};
  frameBuffer_4_78 = _RAND_606[7:0];
  _RAND_607 = {1{`RANDOM}};
  frameBuffer_4_79 = _RAND_607[7:0];
  _RAND_608 = {1{`RANDOM}};
  frameBuffer_4_80 = _RAND_608[7:0];
  _RAND_609 = {1{`RANDOM}};
  frameBuffer_4_81 = _RAND_609[7:0];
  _RAND_610 = {1{`RANDOM}};
  frameBuffer_4_82 = _RAND_610[7:0];
  _RAND_611 = {1{`RANDOM}};
  frameBuffer_4_83 = _RAND_611[7:0];
  _RAND_612 = {1{`RANDOM}};
  frameBuffer_4_84 = _RAND_612[7:0];
  _RAND_613 = {1{`RANDOM}};
  frameBuffer_4_85 = _RAND_613[7:0];
  _RAND_614 = {1{`RANDOM}};
  frameBuffer_4_86 = _RAND_614[7:0];
  _RAND_615 = {1{`RANDOM}};
  frameBuffer_4_87 = _RAND_615[7:0];
  _RAND_616 = {1{`RANDOM}};
  frameBuffer_4_88 = _RAND_616[7:0];
  _RAND_617 = {1{`RANDOM}};
  frameBuffer_4_89 = _RAND_617[7:0];
  _RAND_618 = {1{`RANDOM}};
  frameBuffer_4_90 = _RAND_618[7:0];
  _RAND_619 = {1{`RANDOM}};
  frameBuffer_4_91 = _RAND_619[7:0];
  _RAND_620 = {1{`RANDOM}};
  frameBuffer_4_92 = _RAND_620[7:0];
  _RAND_621 = {1{`RANDOM}};
  frameBuffer_4_93 = _RAND_621[7:0];
  _RAND_622 = {1{`RANDOM}};
  frameBuffer_4_94 = _RAND_622[7:0];
  _RAND_623 = {1{`RANDOM}};
  frameBuffer_4_95 = _RAND_623[7:0];
  _RAND_624 = {1{`RANDOM}};
  frameBuffer_4_96 = _RAND_624[7:0];
  _RAND_625 = {1{`RANDOM}};
  frameBuffer_4_97 = _RAND_625[7:0];
  _RAND_626 = {1{`RANDOM}};
  frameBuffer_4_98 = _RAND_626[7:0];
  _RAND_627 = {1{`RANDOM}};
  frameBuffer_4_99 = _RAND_627[7:0];
  _RAND_628 = {1{`RANDOM}};
  frameBuffer_4_100 = _RAND_628[7:0];
  _RAND_629 = {1{`RANDOM}};
  frameBuffer_4_101 = _RAND_629[7:0];
  _RAND_630 = {1{`RANDOM}};
  frameBuffer_4_102 = _RAND_630[7:0];
  _RAND_631 = {1{`RANDOM}};
  frameBuffer_4_103 = _RAND_631[7:0];
  _RAND_632 = {1{`RANDOM}};
  frameBuffer_4_104 = _RAND_632[7:0];
  _RAND_633 = {1{`RANDOM}};
  frameBuffer_4_105 = _RAND_633[7:0];
  _RAND_634 = {1{`RANDOM}};
  frameBuffer_4_106 = _RAND_634[7:0];
  _RAND_635 = {1{`RANDOM}};
  frameBuffer_4_107 = _RAND_635[7:0];
  _RAND_636 = {1{`RANDOM}};
  frameBuffer_4_108 = _RAND_636[7:0];
  _RAND_637 = {1{`RANDOM}};
  frameBuffer_4_109 = _RAND_637[7:0];
  _RAND_638 = {1{`RANDOM}};
  frameBuffer_4_110 = _RAND_638[7:0];
  _RAND_639 = {1{`RANDOM}};
  frameBuffer_4_111 = _RAND_639[7:0];
  _RAND_640 = {1{`RANDOM}};
  frameBuffer_4_112 = _RAND_640[7:0];
  _RAND_641 = {1{`RANDOM}};
  frameBuffer_4_113 = _RAND_641[7:0];
  _RAND_642 = {1{`RANDOM}};
  frameBuffer_4_114 = _RAND_642[7:0];
  _RAND_643 = {1{`RANDOM}};
  frameBuffer_4_115 = _RAND_643[7:0];
  _RAND_644 = {1{`RANDOM}};
  frameBuffer_4_116 = _RAND_644[7:0];
  _RAND_645 = {1{`RANDOM}};
  frameBuffer_4_117 = _RAND_645[7:0];
  _RAND_646 = {1{`RANDOM}};
  frameBuffer_4_118 = _RAND_646[7:0];
  _RAND_647 = {1{`RANDOM}};
  frameBuffer_4_119 = _RAND_647[7:0];
  _RAND_648 = {1{`RANDOM}};
  frameBuffer_4_120 = _RAND_648[7:0];
  _RAND_649 = {1{`RANDOM}};
  frameBuffer_4_121 = _RAND_649[7:0];
  _RAND_650 = {1{`RANDOM}};
  frameBuffer_4_122 = _RAND_650[7:0];
  _RAND_651 = {1{`RANDOM}};
  frameBuffer_4_123 = _RAND_651[7:0];
  _RAND_652 = {1{`RANDOM}};
  frameBuffer_4_124 = _RAND_652[7:0];
  _RAND_653 = {1{`RANDOM}};
  frameBuffer_4_125 = _RAND_653[7:0];
  _RAND_654 = {1{`RANDOM}};
  frameBuffer_4_126 = _RAND_654[7:0];
  _RAND_655 = {1{`RANDOM}};
  frameBuffer_4_127 = _RAND_655[7:0];
  _RAND_656 = {1{`RANDOM}};
  frameBuffer_5_0 = _RAND_656[7:0];
  _RAND_657 = {1{`RANDOM}};
  frameBuffer_5_1 = _RAND_657[7:0];
  _RAND_658 = {1{`RANDOM}};
  frameBuffer_5_2 = _RAND_658[7:0];
  _RAND_659 = {1{`RANDOM}};
  frameBuffer_5_3 = _RAND_659[7:0];
  _RAND_660 = {1{`RANDOM}};
  frameBuffer_5_4 = _RAND_660[7:0];
  _RAND_661 = {1{`RANDOM}};
  frameBuffer_5_5 = _RAND_661[7:0];
  _RAND_662 = {1{`RANDOM}};
  frameBuffer_5_6 = _RAND_662[7:0];
  _RAND_663 = {1{`RANDOM}};
  frameBuffer_5_7 = _RAND_663[7:0];
  _RAND_664 = {1{`RANDOM}};
  frameBuffer_5_8 = _RAND_664[7:0];
  _RAND_665 = {1{`RANDOM}};
  frameBuffer_5_9 = _RAND_665[7:0];
  _RAND_666 = {1{`RANDOM}};
  frameBuffer_5_10 = _RAND_666[7:0];
  _RAND_667 = {1{`RANDOM}};
  frameBuffer_5_11 = _RAND_667[7:0];
  _RAND_668 = {1{`RANDOM}};
  frameBuffer_5_12 = _RAND_668[7:0];
  _RAND_669 = {1{`RANDOM}};
  frameBuffer_5_13 = _RAND_669[7:0];
  _RAND_670 = {1{`RANDOM}};
  frameBuffer_5_14 = _RAND_670[7:0];
  _RAND_671 = {1{`RANDOM}};
  frameBuffer_5_15 = _RAND_671[7:0];
  _RAND_672 = {1{`RANDOM}};
  frameBuffer_5_16 = _RAND_672[7:0];
  _RAND_673 = {1{`RANDOM}};
  frameBuffer_5_17 = _RAND_673[7:0];
  _RAND_674 = {1{`RANDOM}};
  frameBuffer_5_18 = _RAND_674[7:0];
  _RAND_675 = {1{`RANDOM}};
  frameBuffer_5_19 = _RAND_675[7:0];
  _RAND_676 = {1{`RANDOM}};
  frameBuffer_5_20 = _RAND_676[7:0];
  _RAND_677 = {1{`RANDOM}};
  frameBuffer_5_21 = _RAND_677[7:0];
  _RAND_678 = {1{`RANDOM}};
  frameBuffer_5_22 = _RAND_678[7:0];
  _RAND_679 = {1{`RANDOM}};
  frameBuffer_5_23 = _RAND_679[7:0];
  _RAND_680 = {1{`RANDOM}};
  frameBuffer_5_24 = _RAND_680[7:0];
  _RAND_681 = {1{`RANDOM}};
  frameBuffer_5_25 = _RAND_681[7:0];
  _RAND_682 = {1{`RANDOM}};
  frameBuffer_5_26 = _RAND_682[7:0];
  _RAND_683 = {1{`RANDOM}};
  frameBuffer_5_27 = _RAND_683[7:0];
  _RAND_684 = {1{`RANDOM}};
  frameBuffer_5_28 = _RAND_684[7:0];
  _RAND_685 = {1{`RANDOM}};
  frameBuffer_5_29 = _RAND_685[7:0];
  _RAND_686 = {1{`RANDOM}};
  frameBuffer_5_30 = _RAND_686[7:0];
  _RAND_687 = {1{`RANDOM}};
  frameBuffer_5_31 = _RAND_687[7:0];
  _RAND_688 = {1{`RANDOM}};
  frameBuffer_5_32 = _RAND_688[7:0];
  _RAND_689 = {1{`RANDOM}};
  frameBuffer_5_33 = _RAND_689[7:0];
  _RAND_690 = {1{`RANDOM}};
  frameBuffer_5_34 = _RAND_690[7:0];
  _RAND_691 = {1{`RANDOM}};
  frameBuffer_5_35 = _RAND_691[7:0];
  _RAND_692 = {1{`RANDOM}};
  frameBuffer_5_36 = _RAND_692[7:0];
  _RAND_693 = {1{`RANDOM}};
  frameBuffer_5_37 = _RAND_693[7:0];
  _RAND_694 = {1{`RANDOM}};
  frameBuffer_5_38 = _RAND_694[7:0];
  _RAND_695 = {1{`RANDOM}};
  frameBuffer_5_39 = _RAND_695[7:0];
  _RAND_696 = {1{`RANDOM}};
  frameBuffer_5_40 = _RAND_696[7:0];
  _RAND_697 = {1{`RANDOM}};
  frameBuffer_5_41 = _RAND_697[7:0];
  _RAND_698 = {1{`RANDOM}};
  frameBuffer_5_42 = _RAND_698[7:0];
  _RAND_699 = {1{`RANDOM}};
  frameBuffer_5_43 = _RAND_699[7:0];
  _RAND_700 = {1{`RANDOM}};
  frameBuffer_5_44 = _RAND_700[7:0];
  _RAND_701 = {1{`RANDOM}};
  frameBuffer_5_45 = _RAND_701[7:0];
  _RAND_702 = {1{`RANDOM}};
  frameBuffer_5_46 = _RAND_702[7:0];
  _RAND_703 = {1{`RANDOM}};
  frameBuffer_5_47 = _RAND_703[7:0];
  _RAND_704 = {1{`RANDOM}};
  frameBuffer_5_48 = _RAND_704[7:0];
  _RAND_705 = {1{`RANDOM}};
  frameBuffer_5_49 = _RAND_705[7:0];
  _RAND_706 = {1{`RANDOM}};
  frameBuffer_5_50 = _RAND_706[7:0];
  _RAND_707 = {1{`RANDOM}};
  frameBuffer_5_51 = _RAND_707[7:0];
  _RAND_708 = {1{`RANDOM}};
  frameBuffer_5_52 = _RAND_708[7:0];
  _RAND_709 = {1{`RANDOM}};
  frameBuffer_5_53 = _RAND_709[7:0];
  _RAND_710 = {1{`RANDOM}};
  frameBuffer_5_54 = _RAND_710[7:0];
  _RAND_711 = {1{`RANDOM}};
  frameBuffer_5_55 = _RAND_711[7:0];
  _RAND_712 = {1{`RANDOM}};
  frameBuffer_5_56 = _RAND_712[7:0];
  _RAND_713 = {1{`RANDOM}};
  frameBuffer_5_57 = _RAND_713[7:0];
  _RAND_714 = {1{`RANDOM}};
  frameBuffer_5_58 = _RAND_714[7:0];
  _RAND_715 = {1{`RANDOM}};
  frameBuffer_5_59 = _RAND_715[7:0];
  _RAND_716 = {1{`RANDOM}};
  frameBuffer_5_60 = _RAND_716[7:0];
  _RAND_717 = {1{`RANDOM}};
  frameBuffer_5_61 = _RAND_717[7:0];
  _RAND_718 = {1{`RANDOM}};
  frameBuffer_5_62 = _RAND_718[7:0];
  _RAND_719 = {1{`RANDOM}};
  frameBuffer_5_63 = _RAND_719[7:0];
  _RAND_720 = {1{`RANDOM}};
  frameBuffer_5_64 = _RAND_720[7:0];
  _RAND_721 = {1{`RANDOM}};
  frameBuffer_5_65 = _RAND_721[7:0];
  _RAND_722 = {1{`RANDOM}};
  frameBuffer_5_66 = _RAND_722[7:0];
  _RAND_723 = {1{`RANDOM}};
  frameBuffer_5_67 = _RAND_723[7:0];
  _RAND_724 = {1{`RANDOM}};
  frameBuffer_5_68 = _RAND_724[7:0];
  _RAND_725 = {1{`RANDOM}};
  frameBuffer_5_69 = _RAND_725[7:0];
  _RAND_726 = {1{`RANDOM}};
  frameBuffer_5_70 = _RAND_726[7:0];
  _RAND_727 = {1{`RANDOM}};
  frameBuffer_5_71 = _RAND_727[7:0];
  _RAND_728 = {1{`RANDOM}};
  frameBuffer_5_72 = _RAND_728[7:0];
  _RAND_729 = {1{`RANDOM}};
  frameBuffer_5_73 = _RAND_729[7:0];
  _RAND_730 = {1{`RANDOM}};
  frameBuffer_5_74 = _RAND_730[7:0];
  _RAND_731 = {1{`RANDOM}};
  frameBuffer_5_75 = _RAND_731[7:0];
  _RAND_732 = {1{`RANDOM}};
  frameBuffer_5_76 = _RAND_732[7:0];
  _RAND_733 = {1{`RANDOM}};
  frameBuffer_5_77 = _RAND_733[7:0];
  _RAND_734 = {1{`RANDOM}};
  frameBuffer_5_78 = _RAND_734[7:0];
  _RAND_735 = {1{`RANDOM}};
  frameBuffer_5_79 = _RAND_735[7:0];
  _RAND_736 = {1{`RANDOM}};
  frameBuffer_5_80 = _RAND_736[7:0];
  _RAND_737 = {1{`RANDOM}};
  frameBuffer_5_81 = _RAND_737[7:0];
  _RAND_738 = {1{`RANDOM}};
  frameBuffer_5_82 = _RAND_738[7:0];
  _RAND_739 = {1{`RANDOM}};
  frameBuffer_5_83 = _RAND_739[7:0];
  _RAND_740 = {1{`RANDOM}};
  frameBuffer_5_84 = _RAND_740[7:0];
  _RAND_741 = {1{`RANDOM}};
  frameBuffer_5_85 = _RAND_741[7:0];
  _RAND_742 = {1{`RANDOM}};
  frameBuffer_5_86 = _RAND_742[7:0];
  _RAND_743 = {1{`RANDOM}};
  frameBuffer_5_87 = _RAND_743[7:0];
  _RAND_744 = {1{`RANDOM}};
  frameBuffer_5_88 = _RAND_744[7:0];
  _RAND_745 = {1{`RANDOM}};
  frameBuffer_5_89 = _RAND_745[7:0];
  _RAND_746 = {1{`RANDOM}};
  frameBuffer_5_90 = _RAND_746[7:0];
  _RAND_747 = {1{`RANDOM}};
  frameBuffer_5_91 = _RAND_747[7:0];
  _RAND_748 = {1{`RANDOM}};
  frameBuffer_5_92 = _RAND_748[7:0];
  _RAND_749 = {1{`RANDOM}};
  frameBuffer_5_93 = _RAND_749[7:0];
  _RAND_750 = {1{`RANDOM}};
  frameBuffer_5_94 = _RAND_750[7:0];
  _RAND_751 = {1{`RANDOM}};
  frameBuffer_5_95 = _RAND_751[7:0];
  _RAND_752 = {1{`RANDOM}};
  frameBuffer_5_96 = _RAND_752[7:0];
  _RAND_753 = {1{`RANDOM}};
  frameBuffer_5_97 = _RAND_753[7:0];
  _RAND_754 = {1{`RANDOM}};
  frameBuffer_5_98 = _RAND_754[7:0];
  _RAND_755 = {1{`RANDOM}};
  frameBuffer_5_99 = _RAND_755[7:0];
  _RAND_756 = {1{`RANDOM}};
  frameBuffer_5_100 = _RAND_756[7:0];
  _RAND_757 = {1{`RANDOM}};
  frameBuffer_5_101 = _RAND_757[7:0];
  _RAND_758 = {1{`RANDOM}};
  frameBuffer_5_102 = _RAND_758[7:0];
  _RAND_759 = {1{`RANDOM}};
  frameBuffer_5_103 = _RAND_759[7:0];
  _RAND_760 = {1{`RANDOM}};
  frameBuffer_5_104 = _RAND_760[7:0];
  _RAND_761 = {1{`RANDOM}};
  frameBuffer_5_105 = _RAND_761[7:0];
  _RAND_762 = {1{`RANDOM}};
  frameBuffer_5_106 = _RAND_762[7:0];
  _RAND_763 = {1{`RANDOM}};
  frameBuffer_5_107 = _RAND_763[7:0];
  _RAND_764 = {1{`RANDOM}};
  frameBuffer_5_108 = _RAND_764[7:0];
  _RAND_765 = {1{`RANDOM}};
  frameBuffer_5_109 = _RAND_765[7:0];
  _RAND_766 = {1{`RANDOM}};
  frameBuffer_5_110 = _RAND_766[7:0];
  _RAND_767 = {1{`RANDOM}};
  frameBuffer_5_111 = _RAND_767[7:0];
  _RAND_768 = {1{`RANDOM}};
  frameBuffer_5_112 = _RAND_768[7:0];
  _RAND_769 = {1{`RANDOM}};
  frameBuffer_5_113 = _RAND_769[7:0];
  _RAND_770 = {1{`RANDOM}};
  frameBuffer_5_114 = _RAND_770[7:0];
  _RAND_771 = {1{`RANDOM}};
  frameBuffer_5_115 = _RAND_771[7:0];
  _RAND_772 = {1{`RANDOM}};
  frameBuffer_5_116 = _RAND_772[7:0];
  _RAND_773 = {1{`RANDOM}};
  frameBuffer_5_117 = _RAND_773[7:0];
  _RAND_774 = {1{`RANDOM}};
  frameBuffer_5_118 = _RAND_774[7:0];
  _RAND_775 = {1{`RANDOM}};
  frameBuffer_5_119 = _RAND_775[7:0];
  _RAND_776 = {1{`RANDOM}};
  frameBuffer_5_120 = _RAND_776[7:0];
  _RAND_777 = {1{`RANDOM}};
  frameBuffer_5_121 = _RAND_777[7:0];
  _RAND_778 = {1{`RANDOM}};
  frameBuffer_5_122 = _RAND_778[7:0];
  _RAND_779 = {1{`RANDOM}};
  frameBuffer_5_123 = _RAND_779[7:0];
  _RAND_780 = {1{`RANDOM}};
  frameBuffer_5_124 = _RAND_780[7:0];
  _RAND_781 = {1{`RANDOM}};
  frameBuffer_5_125 = _RAND_781[7:0];
  _RAND_782 = {1{`RANDOM}};
  frameBuffer_5_126 = _RAND_782[7:0];
  _RAND_783 = {1{`RANDOM}};
  frameBuffer_5_127 = _RAND_783[7:0];
  _RAND_784 = {1{`RANDOM}};
  frameBuffer_6_0 = _RAND_784[7:0];
  _RAND_785 = {1{`RANDOM}};
  frameBuffer_6_1 = _RAND_785[7:0];
  _RAND_786 = {1{`RANDOM}};
  frameBuffer_6_2 = _RAND_786[7:0];
  _RAND_787 = {1{`RANDOM}};
  frameBuffer_6_3 = _RAND_787[7:0];
  _RAND_788 = {1{`RANDOM}};
  frameBuffer_6_4 = _RAND_788[7:0];
  _RAND_789 = {1{`RANDOM}};
  frameBuffer_6_5 = _RAND_789[7:0];
  _RAND_790 = {1{`RANDOM}};
  frameBuffer_6_6 = _RAND_790[7:0];
  _RAND_791 = {1{`RANDOM}};
  frameBuffer_6_7 = _RAND_791[7:0];
  _RAND_792 = {1{`RANDOM}};
  frameBuffer_6_8 = _RAND_792[7:0];
  _RAND_793 = {1{`RANDOM}};
  frameBuffer_6_9 = _RAND_793[7:0];
  _RAND_794 = {1{`RANDOM}};
  frameBuffer_6_10 = _RAND_794[7:0];
  _RAND_795 = {1{`RANDOM}};
  frameBuffer_6_11 = _RAND_795[7:0];
  _RAND_796 = {1{`RANDOM}};
  frameBuffer_6_12 = _RAND_796[7:0];
  _RAND_797 = {1{`RANDOM}};
  frameBuffer_6_13 = _RAND_797[7:0];
  _RAND_798 = {1{`RANDOM}};
  frameBuffer_6_14 = _RAND_798[7:0];
  _RAND_799 = {1{`RANDOM}};
  frameBuffer_6_15 = _RAND_799[7:0];
  _RAND_800 = {1{`RANDOM}};
  frameBuffer_6_16 = _RAND_800[7:0];
  _RAND_801 = {1{`RANDOM}};
  frameBuffer_6_17 = _RAND_801[7:0];
  _RAND_802 = {1{`RANDOM}};
  frameBuffer_6_18 = _RAND_802[7:0];
  _RAND_803 = {1{`RANDOM}};
  frameBuffer_6_19 = _RAND_803[7:0];
  _RAND_804 = {1{`RANDOM}};
  frameBuffer_6_20 = _RAND_804[7:0];
  _RAND_805 = {1{`RANDOM}};
  frameBuffer_6_21 = _RAND_805[7:0];
  _RAND_806 = {1{`RANDOM}};
  frameBuffer_6_22 = _RAND_806[7:0];
  _RAND_807 = {1{`RANDOM}};
  frameBuffer_6_23 = _RAND_807[7:0];
  _RAND_808 = {1{`RANDOM}};
  frameBuffer_6_24 = _RAND_808[7:0];
  _RAND_809 = {1{`RANDOM}};
  frameBuffer_6_25 = _RAND_809[7:0];
  _RAND_810 = {1{`RANDOM}};
  frameBuffer_6_26 = _RAND_810[7:0];
  _RAND_811 = {1{`RANDOM}};
  frameBuffer_6_27 = _RAND_811[7:0];
  _RAND_812 = {1{`RANDOM}};
  frameBuffer_6_28 = _RAND_812[7:0];
  _RAND_813 = {1{`RANDOM}};
  frameBuffer_6_29 = _RAND_813[7:0];
  _RAND_814 = {1{`RANDOM}};
  frameBuffer_6_30 = _RAND_814[7:0];
  _RAND_815 = {1{`RANDOM}};
  frameBuffer_6_31 = _RAND_815[7:0];
  _RAND_816 = {1{`RANDOM}};
  frameBuffer_6_32 = _RAND_816[7:0];
  _RAND_817 = {1{`RANDOM}};
  frameBuffer_6_33 = _RAND_817[7:0];
  _RAND_818 = {1{`RANDOM}};
  frameBuffer_6_34 = _RAND_818[7:0];
  _RAND_819 = {1{`RANDOM}};
  frameBuffer_6_35 = _RAND_819[7:0];
  _RAND_820 = {1{`RANDOM}};
  frameBuffer_6_36 = _RAND_820[7:0];
  _RAND_821 = {1{`RANDOM}};
  frameBuffer_6_37 = _RAND_821[7:0];
  _RAND_822 = {1{`RANDOM}};
  frameBuffer_6_38 = _RAND_822[7:0];
  _RAND_823 = {1{`RANDOM}};
  frameBuffer_6_39 = _RAND_823[7:0];
  _RAND_824 = {1{`RANDOM}};
  frameBuffer_6_40 = _RAND_824[7:0];
  _RAND_825 = {1{`RANDOM}};
  frameBuffer_6_41 = _RAND_825[7:0];
  _RAND_826 = {1{`RANDOM}};
  frameBuffer_6_42 = _RAND_826[7:0];
  _RAND_827 = {1{`RANDOM}};
  frameBuffer_6_43 = _RAND_827[7:0];
  _RAND_828 = {1{`RANDOM}};
  frameBuffer_6_44 = _RAND_828[7:0];
  _RAND_829 = {1{`RANDOM}};
  frameBuffer_6_45 = _RAND_829[7:0];
  _RAND_830 = {1{`RANDOM}};
  frameBuffer_6_46 = _RAND_830[7:0];
  _RAND_831 = {1{`RANDOM}};
  frameBuffer_6_47 = _RAND_831[7:0];
  _RAND_832 = {1{`RANDOM}};
  frameBuffer_6_48 = _RAND_832[7:0];
  _RAND_833 = {1{`RANDOM}};
  frameBuffer_6_49 = _RAND_833[7:0];
  _RAND_834 = {1{`RANDOM}};
  frameBuffer_6_50 = _RAND_834[7:0];
  _RAND_835 = {1{`RANDOM}};
  frameBuffer_6_51 = _RAND_835[7:0];
  _RAND_836 = {1{`RANDOM}};
  frameBuffer_6_52 = _RAND_836[7:0];
  _RAND_837 = {1{`RANDOM}};
  frameBuffer_6_53 = _RAND_837[7:0];
  _RAND_838 = {1{`RANDOM}};
  frameBuffer_6_54 = _RAND_838[7:0];
  _RAND_839 = {1{`RANDOM}};
  frameBuffer_6_55 = _RAND_839[7:0];
  _RAND_840 = {1{`RANDOM}};
  frameBuffer_6_56 = _RAND_840[7:0];
  _RAND_841 = {1{`RANDOM}};
  frameBuffer_6_57 = _RAND_841[7:0];
  _RAND_842 = {1{`RANDOM}};
  frameBuffer_6_58 = _RAND_842[7:0];
  _RAND_843 = {1{`RANDOM}};
  frameBuffer_6_59 = _RAND_843[7:0];
  _RAND_844 = {1{`RANDOM}};
  frameBuffer_6_60 = _RAND_844[7:0];
  _RAND_845 = {1{`RANDOM}};
  frameBuffer_6_61 = _RAND_845[7:0];
  _RAND_846 = {1{`RANDOM}};
  frameBuffer_6_62 = _RAND_846[7:0];
  _RAND_847 = {1{`RANDOM}};
  frameBuffer_6_63 = _RAND_847[7:0];
  _RAND_848 = {1{`RANDOM}};
  frameBuffer_6_64 = _RAND_848[7:0];
  _RAND_849 = {1{`RANDOM}};
  frameBuffer_6_65 = _RAND_849[7:0];
  _RAND_850 = {1{`RANDOM}};
  frameBuffer_6_66 = _RAND_850[7:0];
  _RAND_851 = {1{`RANDOM}};
  frameBuffer_6_67 = _RAND_851[7:0];
  _RAND_852 = {1{`RANDOM}};
  frameBuffer_6_68 = _RAND_852[7:0];
  _RAND_853 = {1{`RANDOM}};
  frameBuffer_6_69 = _RAND_853[7:0];
  _RAND_854 = {1{`RANDOM}};
  frameBuffer_6_70 = _RAND_854[7:0];
  _RAND_855 = {1{`RANDOM}};
  frameBuffer_6_71 = _RAND_855[7:0];
  _RAND_856 = {1{`RANDOM}};
  frameBuffer_6_72 = _RAND_856[7:0];
  _RAND_857 = {1{`RANDOM}};
  frameBuffer_6_73 = _RAND_857[7:0];
  _RAND_858 = {1{`RANDOM}};
  frameBuffer_6_74 = _RAND_858[7:0];
  _RAND_859 = {1{`RANDOM}};
  frameBuffer_6_75 = _RAND_859[7:0];
  _RAND_860 = {1{`RANDOM}};
  frameBuffer_6_76 = _RAND_860[7:0];
  _RAND_861 = {1{`RANDOM}};
  frameBuffer_6_77 = _RAND_861[7:0];
  _RAND_862 = {1{`RANDOM}};
  frameBuffer_6_78 = _RAND_862[7:0];
  _RAND_863 = {1{`RANDOM}};
  frameBuffer_6_79 = _RAND_863[7:0];
  _RAND_864 = {1{`RANDOM}};
  frameBuffer_6_80 = _RAND_864[7:0];
  _RAND_865 = {1{`RANDOM}};
  frameBuffer_6_81 = _RAND_865[7:0];
  _RAND_866 = {1{`RANDOM}};
  frameBuffer_6_82 = _RAND_866[7:0];
  _RAND_867 = {1{`RANDOM}};
  frameBuffer_6_83 = _RAND_867[7:0];
  _RAND_868 = {1{`RANDOM}};
  frameBuffer_6_84 = _RAND_868[7:0];
  _RAND_869 = {1{`RANDOM}};
  frameBuffer_6_85 = _RAND_869[7:0];
  _RAND_870 = {1{`RANDOM}};
  frameBuffer_6_86 = _RAND_870[7:0];
  _RAND_871 = {1{`RANDOM}};
  frameBuffer_6_87 = _RAND_871[7:0];
  _RAND_872 = {1{`RANDOM}};
  frameBuffer_6_88 = _RAND_872[7:0];
  _RAND_873 = {1{`RANDOM}};
  frameBuffer_6_89 = _RAND_873[7:0];
  _RAND_874 = {1{`RANDOM}};
  frameBuffer_6_90 = _RAND_874[7:0];
  _RAND_875 = {1{`RANDOM}};
  frameBuffer_6_91 = _RAND_875[7:0];
  _RAND_876 = {1{`RANDOM}};
  frameBuffer_6_92 = _RAND_876[7:0];
  _RAND_877 = {1{`RANDOM}};
  frameBuffer_6_93 = _RAND_877[7:0];
  _RAND_878 = {1{`RANDOM}};
  frameBuffer_6_94 = _RAND_878[7:0];
  _RAND_879 = {1{`RANDOM}};
  frameBuffer_6_95 = _RAND_879[7:0];
  _RAND_880 = {1{`RANDOM}};
  frameBuffer_6_96 = _RAND_880[7:0];
  _RAND_881 = {1{`RANDOM}};
  frameBuffer_6_97 = _RAND_881[7:0];
  _RAND_882 = {1{`RANDOM}};
  frameBuffer_6_98 = _RAND_882[7:0];
  _RAND_883 = {1{`RANDOM}};
  frameBuffer_6_99 = _RAND_883[7:0];
  _RAND_884 = {1{`RANDOM}};
  frameBuffer_6_100 = _RAND_884[7:0];
  _RAND_885 = {1{`RANDOM}};
  frameBuffer_6_101 = _RAND_885[7:0];
  _RAND_886 = {1{`RANDOM}};
  frameBuffer_6_102 = _RAND_886[7:0];
  _RAND_887 = {1{`RANDOM}};
  frameBuffer_6_103 = _RAND_887[7:0];
  _RAND_888 = {1{`RANDOM}};
  frameBuffer_6_104 = _RAND_888[7:0];
  _RAND_889 = {1{`RANDOM}};
  frameBuffer_6_105 = _RAND_889[7:0];
  _RAND_890 = {1{`RANDOM}};
  frameBuffer_6_106 = _RAND_890[7:0];
  _RAND_891 = {1{`RANDOM}};
  frameBuffer_6_107 = _RAND_891[7:0];
  _RAND_892 = {1{`RANDOM}};
  frameBuffer_6_108 = _RAND_892[7:0];
  _RAND_893 = {1{`RANDOM}};
  frameBuffer_6_109 = _RAND_893[7:0];
  _RAND_894 = {1{`RANDOM}};
  frameBuffer_6_110 = _RAND_894[7:0];
  _RAND_895 = {1{`RANDOM}};
  frameBuffer_6_111 = _RAND_895[7:0];
  _RAND_896 = {1{`RANDOM}};
  frameBuffer_6_112 = _RAND_896[7:0];
  _RAND_897 = {1{`RANDOM}};
  frameBuffer_6_113 = _RAND_897[7:0];
  _RAND_898 = {1{`RANDOM}};
  frameBuffer_6_114 = _RAND_898[7:0];
  _RAND_899 = {1{`RANDOM}};
  frameBuffer_6_115 = _RAND_899[7:0];
  _RAND_900 = {1{`RANDOM}};
  frameBuffer_6_116 = _RAND_900[7:0];
  _RAND_901 = {1{`RANDOM}};
  frameBuffer_6_117 = _RAND_901[7:0];
  _RAND_902 = {1{`RANDOM}};
  frameBuffer_6_118 = _RAND_902[7:0];
  _RAND_903 = {1{`RANDOM}};
  frameBuffer_6_119 = _RAND_903[7:0];
  _RAND_904 = {1{`RANDOM}};
  frameBuffer_6_120 = _RAND_904[7:0];
  _RAND_905 = {1{`RANDOM}};
  frameBuffer_6_121 = _RAND_905[7:0];
  _RAND_906 = {1{`RANDOM}};
  frameBuffer_6_122 = _RAND_906[7:0];
  _RAND_907 = {1{`RANDOM}};
  frameBuffer_6_123 = _RAND_907[7:0];
  _RAND_908 = {1{`RANDOM}};
  frameBuffer_6_124 = _RAND_908[7:0];
  _RAND_909 = {1{`RANDOM}};
  frameBuffer_6_125 = _RAND_909[7:0];
  _RAND_910 = {1{`RANDOM}};
  frameBuffer_6_126 = _RAND_910[7:0];
  _RAND_911 = {1{`RANDOM}};
  frameBuffer_6_127 = _RAND_911[7:0];
  _RAND_912 = {1{`RANDOM}};
  frameBuffer_7_0 = _RAND_912[7:0];
  _RAND_913 = {1{`RANDOM}};
  frameBuffer_7_1 = _RAND_913[7:0];
  _RAND_914 = {1{`RANDOM}};
  frameBuffer_7_2 = _RAND_914[7:0];
  _RAND_915 = {1{`RANDOM}};
  frameBuffer_7_3 = _RAND_915[7:0];
  _RAND_916 = {1{`RANDOM}};
  frameBuffer_7_4 = _RAND_916[7:0];
  _RAND_917 = {1{`RANDOM}};
  frameBuffer_7_5 = _RAND_917[7:0];
  _RAND_918 = {1{`RANDOM}};
  frameBuffer_7_6 = _RAND_918[7:0];
  _RAND_919 = {1{`RANDOM}};
  frameBuffer_7_7 = _RAND_919[7:0];
  _RAND_920 = {1{`RANDOM}};
  frameBuffer_7_8 = _RAND_920[7:0];
  _RAND_921 = {1{`RANDOM}};
  frameBuffer_7_9 = _RAND_921[7:0];
  _RAND_922 = {1{`RANDOM}};
  frameBuffer_7_10 = _RAND_922[7:0];
  _RAND_923 = {1{`RANDOM}};
  frameBuffer_7_11 = _RAND_923[7:0];
  _RAND_924 = {1{`RANDOM}};
  frameBuffer_7_12 = _RAND_924[7:0];
  _RAND_925 = {1{`RANDOM}};
  frameBuffer_7_13 = _RAND_925[7:0];
  _RAND_926 = {1{`RANDOM}};
  frameBuffer_7_14 = _RAND_926[7:0];
  _RAND_927 = {1{`RANDOM}};
  frameBuffer_7_15 = _RAND_927[7:0];
  _RAND_928 = {1{`RANDOM}};
  frameBuffer_7_16 = _RAND_928[7:0];
  _RAND_929 = {1{`RANDOM}};
  frameBuffer_7_17 = _RAND_929[7:0];
  _RAND_930 = {1{`RANDOM}};
  frameBuffer_7_18 = _RAND_930[7:0];
  _RAND_931 = {1{`RANDOM}};
  frameBuffer_7_19 = _RAND_931[7:0];
  _RAND_932 = {1{`RANDOM}};
  frameBuffer_7_20 = _RAND_932[7:0];
  _RAND_933 = {1{`RANDOM}};
  frameBuffer_7_21 = _RAND_933[7:0];
  _RAND_934 = {1{`RANDOM}};
  frameBuffer_7_22 = _RAND_934[7:0];
  _RAND_935 = {1{`RANDOM}};
  frameBuffer_7_23 = _RAND_935[7:0];
  _RAND_936 = {1{`RANDOM}};
  frameBuffer_7_24 = _RAND_936[7:0];
  _RAND_937 = {1{`RANDOM}};
  frameBuffer_7_25 = _RAND_937[7:0];
  _RAND_938 = {1{`RANDOM}};
  frameBuffer_7_26 = _RAND_938[7:0];
  _RAND_939 = {1{`RANDOM}};
  frameBuffer_7_27 = _RAND_939[7:0];
  _RAND_940 = {1{`RANDOM}};
  frameBuffer_7_28 = _RAND_940[7:0];
  _RAND_941 = {1{`RANDOM}};
  frameBuffer_7_29 = _RAND_941[7:0];
  _RAND_942 = {1{`RANDOM}};
  frameBuffer_7_30 = _RAND_942[7:0];
  _RAND_943 = {1{`RANDOM}};
  frameBuffer_7_31 = _RAND_943[7:0];
  _RAND_944 = {1{`RANDOM}};
  frameBuffer_7_32 = _RAND_944[7:0];
  _RAND_945 = {1{`RANDOM}};
  frameBuffer_7_33 = _RAND_945[7:0];
  _RAND_946 = {1{`RANDOM}};
  frameBuffer_7_34 = _RAND_946[7:0];
  _RAND_947 = {1{`RANDOM}};
  frameBuffer_7_35 = _RAND_947[7:0];
  _RAND_948 = {1{`RANDOM}};
  frameBuffer_7_36 = _RAND_948[7:0];
  _RAND_949 = {1{`RANDOM}};
  frameBuffer_7_37 = _RAND_949[7:0];
  _RAND_950 = {1{`RANDOM}};
  frameBuffer_7_38 = _RAND_950[7:0];
  _RAND_951 = {1{`RANDOM}};
  frameBuffer_7_39 = _RAND_951[7:0];
  _RAND_952 = {1{`RANDOM}};
  frameBuffer_7_40 = _RAND_952[7:0];
  _RAND_953 = {1{`RANDOM}};
  frameBuffer_7_41 = _RAND_953[7:0];
  _RAND_954 = {1{`RANDOM}};
  frameBuffer_7_42 = _RAND_954[7:0];
  _RAND_955 = {1{`RANDOM}};
  frameBuffer_7_43 = _RAND_955[7:0];
  _RAND_956 = {1{`RANDOM}};
  frameBuffer_7_44 = _RAND_956[7:0];
  _RAND_957 = {1{`RANDOM}};
  frameBuffer_7_45 = _RAND_957[7:0];
  _RAND_958 = {1{`RANDOM}};
  frameBuffer_7_46 = _RAND_958[7:0];
  _RAND_959 = {1{`RANDOM}};
  frameBuffer_7_47 = _RAND_959[7:0];
  _RAND_960 = {1{`RANDOM}};
  frameBuffer_7_48 = _RAND_960[7:0];
  _RAND_961 = {1{`RANDOM}};
  frameBuffer_7_49 = _RAND_961[7:0];
  _RAND_962 = {1{`RANDOM}};
  frameBuffer_7_50 = _RAND_962[7:0];
  _RAND_963 = {1{`RANDOM}};
  frameBuffer_7_51 = _RAND_963[7:0];
  _RAND_964 = {1{`RANDOM}};
  frameBuffer_7_52 = _RAND_964[7:0];
  _RAND_965 = {1{`RANDOM}};
  frameBuffer_7_53 = _RAND_965[7:0];
  _RAND_966 = {1{`RANDOM}};
  frameBuffer_7_54 = _RAND_966[7:0];
  _RAND_967 = {1{`RANDOM}};
  frameBuffer_7_55 = _RAND_967[7:0];
  _RAND_968 = {1{`RANDOM}};
  frameBuffer_7_56 = _RAND_968[7:0];
  _RAND_969 = {1{`RANDOM}};
  frameBuffer_7_57 = _RAND_969[7:0];
  _RAND_970 = {1{`RANDOM}};
  frameBuffer_7_58 = _RAND_970[7:0];
  _RAND_971 = {1{`RANDOM}};
  frameBuffer_7_59 = _RAND_971[7:0];
  _RAND_972 = {1{`RANDOM}};
  frameBuffer_7_60 = _RAND_972[7:0];
  _RAND_973 = {1{`RANDOM}};
  frameBuffer_7_61 = _RAND_973[7:0];
  _RAND_974 = {1{`RANDOM}};
  frameBuffer_7_62 = _RAND_974[7:0];
  _RAND_975 = {1{`RANDOM}};
  frameBuffer_7_63 = _RAND_975[7:0];
  _RAND_976 = {1{`RANDOM}};
  frameBuffer_7_64 = _RAND_976[7:0];
  _RAND_977 = {1{`RANDOM}};
  frameBuffer_7_65 = _RAND_977[7:0];
  _RAND_978 = {1{`RANDOM}};
  frameBuffer_7_66 = _RAND_978[7:0];
  _RAND_979 = {1{`RANDOM}};
  frameBuffer_7_67 = _RAND_979[7:0];
  _RAND_980 = {1{`RANDOM}};
  frameBuffer_7_68 = _RAND_980[7:0];
  _RAND_981 = {1{`RANDOM}};
  frameBuffer_7_69 = _RAND_981[7:0];
  _RAND_982 = {1{`RANDOM}};
  frameBuffer_7_70 = _RAND_982[7:0];
  _RAND_983 = {1{`RANDOM}};
  frameBuffer_7_71 = _RAND_983[7:0];
  _RAND_984 = {1{`RANDOM}};
  frameBuffer_7_72 = _RAND_984[7:0];
  _RAND_985 = {1{`RANDOM}};
  frameBuffer_7_73 = _RAND_985[7:0];
  _RAND_986 = {1{`RANDOM}};
  frameBuffer_7_74 = _RAND_986[7:0];
  _RAND_987 = {1{`RANDOM}};
  frameBuffer_7_75 = _RAND_987[7:0];
  _RAND_988 = {1{`RANDOM}};
  frameBuffer_7_76 = _RAND_988[7:0];
  _RAND_989 = {1{`RANDOM}};
  frameBuffer_7_77 = _RAND_989[7:0];
  _RAND_990 = {1{`RANDOM}};
  frameBuffer_7_78 = _RAND_990[7:0];
  _RAND_991 = {1{`RANDOM}};
  frameBuffer_7_79 = _RAND_991[7:0];
  _RAND_992 = {1{`RANDOM}};
  frameBuffer_7_80 = _RAND_992[7:0];
  _RAND_993 = {1{`RANDOM}};
  frameBuffer_7_81 = _RAND_993[7:0];
  _RAND_994 = {1{`RANDOM}};
  frameBuffer_7_82 = _RAND_994[7:0];
  _RAND_995 = {1{`RANDOM}};
  frameBuffer_7_83 = _RAND_995[7:0];
  _RAND_996 = {1{`RANDOM}};
  frameBuffer_7_84 = _RAND_996[7:0];
  _RAND_997 = {1{`RANDOM}};
  frameBuffer_7_85 = _RAND_997[7:0];
  _RAND_998 = {1{`RANDOM}};
  frameBuffer_7_86 = _RAND_998[7:0];
  _RAND_999 = {1{`RANDOM}};
  frameBuffer_7_87 = _RAND_999[7:0];
  _RAND_1000 = {1{`RANDOM}};
  frameBuffer_7_88 = _RAND_1000[7:0];
  _RAND_1001 = {1{`RANDOM}};
  frameBuffer_7_89 = _RAND_1001[7:0];
  _RAND_1002 = {1{`RANDOM}};
  frameBuffer_7_90 = _RAND_1002[7:0];
  _RAND_1003 = {1{`RANDOM}};
  frameBuffer_7_91 = _RAND_1003[7:0];
  _RAND_1004 = {1{`RANDOM}};
  frameBuffer_7_92 = _RAND_1004[7:0];
  _RAND_1005 = {1{`RANDOM}};
  frameBuffer_7_93 = _RAND_1005[7:0];
  _RAND_1006 = {1{`RANDOM}};
  frameBuffer_7_94 = _RAND_1006[7:0];
  _RAND_1007 = {1{`RANDOM}};
  frameBuffer_7_95 = _RAND_1007[7:0];
  _RAND_1008 = {1{`RANDOM}};
  frameBuffer_7_96 = _RAND_1008[7:0];
  _RAND_1009 = {1{`RANDOM}};
  frameBuffer_7_97 = _RAND_1009[7:0];
  _RAND_1010 = {1{`RANDOM}};
  frameBuffer_7_98 = _RAND_1010[7:0];
  _RAND_1011 = {1{`RANDOM}};
  frameBuffer_7_99 = _RAND_1011[7:0];
  _RAND_1012 = {1{`RANDOM}};
  frameBuffer_7_100 = _RAND_1012[7:0];
  _RAND_1013 = {1{`RANDOM}};
  frameBuffer_7_101 = _RAND_1013[7:0];
  _RAND_1014 = {1{`RANDOM}};
  frameBuffer_7_102 = _RAND_1014[7:0];
  _RAND_1015 = {1{`RANDOM}};
  frameBuffer_7_103 = _RAND_1015[7:0];
  _RAND_1016 = {1{`RANDOM}};
  frameBuffer_7_104 = _RAND_1016[7:0];
  _RAND_1017 = {1{`RANDOM}};
  frameBuffer_7_105 = _RAND_1017[7:0];
  _RAND_1018 = {1{`RANDOM}};
  frameBuffer_7_106 = _RAND_1018[7:0];
  _RAND_1019 = {1{`RANDOM}};
  frameBuffer_7_107 = _RAND_1019[7:0];
  _RAND_1020 = {1{`RANDOM}};
  frameBuffer_7_108 = _RAND_1020[7:0];
  _RAND_1021 = {1{`RANDOM}};
  frameBuffer_7_109 = _RAND_1021[7:0];
  _RAND_1022 = {1{`RANDOM}};
  frameBuffer_7_110 = _RAND_1022[7:0];
  _RAND_1023 = {1{`RANDOM}};
  frameBuffer_7_111 = _RAND_1023[7:0];
  _RAND_1024 = {1{`RANDOM}};
  frameBuffer_7_112 = _RAND_1024[7:0];
  _RAND_1025 = {1{`RANDOM}};
  frameBuffer_7_113 = _RAND_1025[7:0];
  _RAND_1026 = {1{`RANDOM}};
  frameBuffer_7_114 = _RAND_1026[7:0];
  _RAND_1027 = {1{`RANDOM}};
  frameBuffer_7_115 = _RAND_1027[7:0];
  _RAND_1028 = {1{`RANDOM}};
  frameBuffer_7_116 = _RAND_1028[7:0];
  _RAND_1029 = {1{`RANDOM}};
  frameBuffer_7_117 = _RAND_1029[7:0];
  _RAND_1030 = {1{`RANDOM}};
  frameBuffer_7_118 = _RAND_1030[7:0];
  _RAND_1031 = {1{`RANDOM}};
  frameBuffer_7_119 = _RAND_1031[7:0];
  _RAND_1032 = {1{`RANDOM}};
  frameBuffer_7_120 = _RAND_1032[7:0];
  _RAND_1033 = {1{`RANDOM}};
  frameBuffer_7_121 = _RAND_1033[7:0];
  _RAND_1034 = {1{`RANDOM}};
  frameBuffer_7_122 = _RAND_1034[7:0];
  _RAND_1035 = {1{`RANDOM}};
  frameBuffer_7_123 = _RAND_1035[7:0];
  _RAND_1036 = {1{`RANDOM}};
  frameBuffer_7_124 = _RAND_1036[7:0];
  _RAND_1037 = {1{`RANDOM}};
  frameBuffer_7_125 = _RAND_1037[7:0];
  _RAND_1038 = {1{`RANDOM}};
  frameBuffer_7_126 = _RAND_1038[7:0];
  _RAND_1039 = {1{`RANDOM}};
  frameBuffer_7_127 = _RAND_1039[7:0];
  _RAND_1040 = {1{`RANDOM}};
  frameBuffer_8_0 = _RAND_1040[7:0];
  _RAND_1041 = {1{`RANDOM}};
  frameBuffer_8_1 = _RAND_1041[7:0];
  _RAND_1042 = {1{`RANDOM}};
  frameBuffer_8_2 = _RAND_1042[7:0];
  _RAND_1043 = {1{`RANDOM}};
  frameBuffer_8_3 = _RAND_1043[7:0];
  _RAND_1044 = {1{`RANDOM}};
  frameBuffer_8_4 = _RAND_1044[7:0];
  _RAND_1045 = {1{`RANDOM}};
  frameBuffer_8_5 = _RAND_1045[7:0];
  _RAND_1046 = {1{`RANDOM}};
  frameBuffer_8_6 = _RAND_1046[7:0];
  _RAND_1047 = {1{`RANDOM}};
  frameBuffer_8_7 = _RAND_1047[7:0];
  _RAND_1048 = {1{`RANDOM}};
  frameBuffer_8_8 = _RAND_1048[7:0];
  _RAND_1049 = {1{`RANDOM}};
  frameBuffer_8_9 = _RAND_1049[7:0];
  _RAND_1050 = {1{`RANDOM}};
  frameBuffer_8_10 = _RAND_1050[7:0];
  _RAND_1051 = {1{`RANDOM}};
  frameBuffer_8_11 = _RAND_1051[7:0];
  _RAND_1052 = {1{`RANDOM}};
  frameBuffer_8_12 = _RAND_1052[7:0];
  _RAND_1053 = {1{`RANDOM}};
  frameBuffer_8_13 = _RAND_1053[7:0];
  _RAND_1054 = {1{`RANDOM}};
  frameBuffer_8_14 = _RAND_1054[7:0];
  _RAND_1055 = {1{`RANDOM}};
  frameBuffer_8_15 = _RAND_1055[7:0];
  _RAND_1056 = {1{`RANDOM}};
  frameBuffer_8_16 = _RAND_1056[7:0];
  _RAND_1057 = {1{`RANDOM}};
  frameBuffer_8_17 = _RAND_1057[7:0];
  _RAND_1058 = {1{`RANDOM}};
  frameBuffer_8_18 = _RAND_1058[7:0];
  _RAND_1059 = {1{`RANDOM}};
  frameBuffer_8_19 = _RAND_1059[7:0];
  _RAND_1060 = {1{`RANDOM}};
  frameBuffer_8_20 = _RAND_1060[7:0];
  _RAND_1061 = {1{`RANDOM}};
  frameBuffer_8_21 = _RAND_1061[7:0];
  _RAND_1062 = {1{`RANDOM}};
  frameBuffer_8_22 = _RAND_1062[7:0];
  _RAND_1063 = {1{`RANDOM}};
  frameBuffer_8_23 = _RAND_1063[7:0];
  _RAND_1064 = {1{`RANDOM}};
  frameBuffer_8_24 = _RAND_1064[7:0];
  _RAND_1065 = {1{`RANDOM}};
  frameBuffer_8_25 = _RAND_1065[7:0];
  _RAND_1066 = {1{`RANDOM}};
  frameBuffer_8_26 = _RAND_1066[7:0];
  _RAND_1067 = {1{`RANDOM}};
  frameBuffer_8_27 = _RAND_1067[7:0];
  _RAND_1068 = {1{`RANDOM}};
  frameBuffer_8_28 = _RAND_1068[7:0];
  _RAND_1069 = {1{`RANDOM}};
  frameBuffer_8_29 = _RAND_1069[7:0];
  _RAND_1070 = {1{`RANDOM}};
  frameBuffer_8_30 = _RAND_1070[7:0];
  _RAND_1071 = {1{`RANDOM}};
  frameBuffer_8_31 = _RAND_1071[7:0];
  _RAND_1072 = {1{`RANDOM}};
  frameBuffer_8_32 = _RAND_1072[7:0];
  _RAND_1073 = {1{`RANDOM}};
  frameBuffer_8_33 = _RAND_1073[7:0];
  _RAND_1074 = {1{`RANDOM}};
  frameBuffer_8_34 = _RAND_1074[7:0];
  _RAND_1075 = {1{`RANDOM}};
  frameBuffer_8_35 = _RAND_1075[7:0];
  _RAND_1076 = {1{`RANDOM}};
  frameBuffer_8_36 = _RAND_1076[7:0];
  _RAND_1077 = {1{`RANDOM}};
  frameBuffer_8_37 = _RAND_1077[7:0];
  _RAND_1078 = {1{`RANDOM}};
  frameBuffer_8_38 = _RAND_1078[7:0];
  _RAND_1079 = {1{`RANDOM}};
  frameBuffer_8_39 = _RAND_1079[7:0];
  _RAND_1080 = {1{`RANDOM}};
  frameBuffer_8_40 = _RAND_1080[7:0];
  _RAND_1081 = {1{`RANDOM}};
  frameBuffer_8_41 = _RAND_1081[7:0];
  _RAND_1082 = {1{`RANDOM}};
  frameBuffer_8_42 = _RAND_1082[7:0];
  _RAND_1083 = {1{`RANDOM}};
  frameBuffer_8_43 = _RAND_1083[7:0];
  _RAND_1084 = {1{`RANDOM}};
  frameBuffer_8_44 = _RAND_1084[7:0];
  _RAND_1085 = {1{`RANDOM}};
  frameBuffer_8_45 = _RAND_1085[7:0];
  _RAND_1086 = {1{`RANDOM}};
  frameBuffer_8_46 = _RAND_1086[7:0];
  _RAND_1087 = {1{`RANDOM}};
  frameBuffer_8_47 = _RAND_1087[7:0];
  _RAND_1088 = {1{`RANDOM}};
  frameBuffer_8_48 = _RAND_1088[7:0];
  _RAND_1089 = {1{`RANDOM}};
  frameBuffer_8_49 = _RAND_1089[7:0];
  _RAND_1090 = {1{`RANDOM}};
  frameBuffer_8_50 = _RAND_1090[7:0];
  _RAND_1091 = {1{`RANDOM}};
  frameBuffer_8_51 = _RAND_1091[7:0];
  _RAND_1092 = {1{`RANDOM}};
  frameBuffer_8_52 = _RAND_1092[7:0];
  _RAND_1093 = {1{`RANDOM}};
  frameBuffer_8_53 = _RAND_1093[7:0];
  _RAND_1094 = {1{`RANDOM}};
  frameBuffer_8_54 = _RAND_1094[7:0];
  _RAND_1095 = {1{`RANDOM}};
  frameBuffer_8_55 = _RAND_1095[7:0];
  _RAND_1096 = {1{`RANDOM}};
  frameBuffer_8_56 = _RAND_1096[7:0];
  _RAND_1097 = {1{`RANDOM}};
  frameBuffer_8_57 = _RAND_1097[7:0];
  _RAND_1098 = {1{`RANDOM}};
  frameBuffer_8_58 = _RAND_1098[7:0];
  _RAND_1099 = {1{`RANDOM}};
  frameBuffer_8_59 = _RAND_1099[7:0];
  _RAND_1100 = {1{`RANDOM}};
  frameBuffer_8_60 = _RAND_1100[7:0];
  _RAND_1101 = {1{`RANDOM}};
  frameBuffer_8_61 = _RAND_1101[7:0];
  _RAND_1102 = {1{`RANDOM}};
  frameBuffer_8_62 = _RAND_1102[7:0];
  _RAND_1103 = {1{`RANDOM}};
  frameBuffer_8_63 = _RAND_1103[7:0];
  _RAND_1104 = {1{`RANDOM}};
  frameBuffer_8_64 = _RAND_1104[7:0];
  _RAND_1105 = {1{`RANDOM}};
  frameBuffer_8_65 = _RAND_1105[7:0];
  _RAND_1106 = {1{`RANDOM}};
  frameBuffer_8_66 = _RAND_1106[7:0];
  _RAND_1107 = {1{`RANDOM}};
  frameBuffer_8_67 = _RAND_1107[7:0];
  _RAND_1108 = {1{`RANDOM}};
  frameBuffer_8_68 = _RAND_1108[7:0];
  _RAND_1109 = {1{`RANDOM}};
  frameBuffer_8_69 = _RAND_1109[7:0];
  _RAND_1110 = {1{`RANDOM}};
  frameBuffer_8_70 = _RAND_1110[7:0];
  _RAND_1111 = {1{`RANDOM}};
  frameBuffer_8_71 = _RAND_1111[7:0];
  _RAND_1112 = {1{`RANDOM}};
  frameBuffer_8_72 = _RAND_1112[7:0];
  _RAND_1113 = {1{`RANDOM}};
  frameBuffer_8_73 = _RAND_1113[7:0];
  _RAND_1114 = {1{`RANDOM}};
  frameBuffer_8_74 = _RAND_1114[7:0];
  _RAND_1115 = {1{`RANDOM}};
  frameBuffer_8_75 = _RAND_1115[7:0];
  _RAND_1116 = {1{`RANDOM}};
  frameBuffer_8_76 = _RAND_1116[7:0];
  _RAND_1117 = {1{`RANDOM}};
  frameBuffer_8_77 = _RAND_1117[7:0];
  _RAND_1118 = {1{`RANDOM}};
  frameBuffer_8_78 = _RAND_1118[7:0];
  _RAND_1119 = {1{`RANDOM}};
  frameBuffer_8_79 = _RAND_1119[7:0];
  _RAND_1120 = {1{`RANDOM}};
  frameBuffer_8_80 = _RAND_1120[7:0];
  _RAND_1121 = {1{`RANDOM}};
  frameBuffer_8_81 = _RAND_1121[7:0];
  _RAND_1122 = {1{`RANDOM}};
  frameBuffer_8_82 = _RAND_1122[7:0];
  _RAND_1123 = {1{`RANDOM}};
  frameBuffer_8_83 = _RAND_1123[7:0];
  _RAND_1124 = {1{`RANDOM}};
  frameBuffer_8_84 = _RAND_1124[7:0];
  _RAND_1125 = {1{`RANDOM}};
  frameBuffer_8_85 = _RAND_1125[7:0];
  _RAND_1126 = {1{`RANDOM}};
  frameBuffer_8_86 = _RAND_1126[7:0];
  _RAND_1127 = {1{`RANDOM}};
  frameBuffer_8_87 = _RAND_1127[7:0];
  _RAND_1128 = {1{`RANDOM}};
  frameBuffer_8_88 = _RAND_1128[7:0];
  _RAND_1129 = {1{`RANDOM}};
  frameBuffer_8_89 = _RAND_1129[7:0];
  _RAND_1130 = {1{`RANDOM}};
  frameBuffer_8_90 = _RAND_1130[7:0];
  _RAND_1131 = {1{`RANDOM}};
  frameBuffer_8_91 = _RAND_1131[7:0];
  _RAND_1132 = {1{`RANDOM}};
  frameBuffer_8_92 = _RAND_1132[7:0];
  _RAND_1133 = {1{`RANDOM}};
  frameBuffer_8_93 = _RAND_1133[7:0];
  _RAND_1134 = {1{`RANDOM}};
  frameBuffer_8_94 = _RAND_1134[7:0];
  _RAND_1135 = {1{`RANDOM}};
  frameBuffer_8_95 = _RAND_1135[7:0];
  _RAND_1136 = {1{`RANDOM}};
  frameBuffer_8_96 = _RAND_1136[7:0];
  _RAND_1137 = {1{`RANDOM}};
  frameBuffer_8_97 = _RAND_1137[7:0];
  _RAND_1138 = {1{`RANDOM}};
  frameBuffer_8_98 = _RAND_1138[7:0];
  _RAND_1139 = {1{`RANDOM}};
  frameBuffer_8_99 = _RAND_1139[7:0];
  _RAND_1140 = {1{`RANDOM}};
  frameBuffer_8_100 = _RAND_1140[7:0];
  _RAND_1141 = {1{`RANDOM}};
  frameBuffer_8_101 = _RAND_1141[7:0];
  _RAND_1142 = {1{`RANDOM}};
  frameBuffer_8_102 = _RAND_1142[7:0];
  _RAND_1143 = {1{`RANDOM}};
  frameBuffer_8_103 = _RAND_1143[7:0];
  _RAND_1144 = {1{`RANDOM}};
  frameBuffer_8_104 = _RAND_1144[7:0];
  _RAND_1145 = {1{`RANDOM}};
  frameBuffer_8_105 = _RAND_1145[7:0];
  _RAND_1146 = {1{`RANDOM}};
  frameBuffer_8_106 = _RAND_1146[7:0];
  _RAND_1147 = {1{`RANDOM}};
  frameBuffer_8_107 = _RAND_1147[7:0];
  _RAND_1148 = {1{`RANDOM}};
  frameBuffer_8_108 = _RAND_1148[7:0];
  _RAND_1149 = {1{`RANDOM}};
  frameBuffer_8_109 = _RAND_1149[7:0];
  _RAND_1150 = {1{`RANDOM}};
  frameBuffer_8_110 = _RAND_1150[7:0];
  _RAND_1151 = {1{`RANDOM}};
  frameBuffer_8_111 = _RAND_1151[7:0];
  _RAND_1152 = {1{`RANDOM}};
  frameBuffer_8_112 = _RAND_1152[7:0];
  _RAND_1153 = {1{`RANDOM}};
  frameBuffer_8_113 = _RAND_1153[7:0];
  _RAND_1154 = {1{`RANDOM}};
  frameBuffer_8_114 = _RAND_1154[7:0];
  _RAND_1155 = {1{`RANDOM}};
  frameBuffer_8_115 = _RAND_1155[7:0];
  _RAND_1156 = {1{`RANDOM}};
  frameBuffer_8_116 = _RAND_1156[7:0];
  _RAND_1157 = {1{`RANDOM}};
  frameBuffer_8_117 = _RAND_1157[7:0];
  _RAND_1158 = {1{`RANDOM}};
  frameBuffer_8_118 = _RAND_1158[7:0];
  _RAND_1159 = {1{`RANDOM}};
  frameBuffer_8_119 = _RAND_1159[7:0];
  _RAND_1160 = {1{`RANDOM}};
  frameBuffer_8_120 = _RAND_1160[7:0];
  _RAND_1161 = {1{`RANDOM}};
  frameBuffer_8_121 = _RAND_1161[7:0];
  _RAND_1162 = {1{`RANDOM}};
  frameBuffer_8_122 = _RAND_1162[7:0];
  _RAND_1163 = {1{`RANDOM}};
  frameBuffer_8_123 = _RAND_1163[7:0];
  _RAND_1164 = {1{`RANDOM}};
  frameBuffer_8_124 = _RAND_1164[7:0];
  _RAND_1165 = {1{`RANDOM}};
  frameBuffer_8_125 = _RAND_1165[7:0];
  _RAND_1166 = {1{`RANDOM}};
  frameBuffer_8_126 = _RAND_1166[7:0];
  _RAND_1167 = {1{`RANDOM}};
  frameBuffer_8_127 = _RAND_1167[7:0];
  _RAND_1168 = {1{`RANDOM}};
  frameBuffer_9_0 = _RAND_1168[7:0];
  _RAND_1169 = {1{`RANDOM}};
  frameBuffer_9_1 = _RAND_1169[7:0];
  _RAND_1170 = {1{`RANDOM}};
  frameBuffer_9_2 = _RAND_1170[7:0];
  _RAND_1171 = {1{`RANDOM}};
  frameBuffer_9_3 = _RAND_1171[7:0];
  _RAND_1172 = {1{`RANDOM}};
  frameBuffer_9_4 = _RAND_1172[7:0];
  _RAND_1173 = {1{`RANDOM}};
  frameBuffer_9_5 = _RAND_1173[7:0];
  _RAND_1174 = {1{`RANDOM}};
  frameBuffer_9_6 = _RAND_1174[7:0];
  _RAND_1175 = {1{`RANDOM}};
  frameBuffer_9_7 = _RAND_1175[7:0];
  _RAND_1176 = {1{`RANDOM}};
  frameBuffer_9_8 = _RAND_1176[7:0];
  _RAND_1177 = {1{`RANDOM}};
  frameBuffer_9_9 = _RAND_1177[7:0];
  _RAND_1178 = {1{`RANDOM}};
  frameBuffer_9_10 = _RAND_1178[7:0];
  _RAND_1179 = {1{`RANDOM}};
  frameBuffer_9_11 = _RAND_1179[7:0];
  _RAND_1180 = {1{`RANDOM}};
  frameBuffer_9_12 = _RAND_1180[7:0];
  _RAND_1181 = {1{`RANDOM}};
  frameBuffer_9_13 = _RAND_1181[7:0];
  _RAND_1182 = {1{`RANDOM}};
  frameBuffer_9_14 = _RAND_1182[7:0];
  _RAND_1183 = {1{`RANDOM}};
  frameBuffer_9_15 = _RAND_1183[7:0];
  _RAND_1184 = {1{`RANDOM}};
  frameBuffer_9_16 = _RAND_1184[7:0];
  _RAND_1185 = {1{`RANDOM}};
  frameBuffer_9_17 = _RAND_1185[7:0];
  _RAND_1186 = {1{`RANDOM}};
  frameBuffer_9_18 = _RAND_1186[7:0];
  _RAND_1187 = {1{`RANDOM}};
  frameBuffer_9_19 = _RAND_1187[7:0];
  _RAND_1188 = {1{`RANDOM}};
  frameBuffer_9_20 = _RAND_1188[7:0];
  _RAND_1189 = {1{`RANDOM}};
  frameBuffer_9_21 = _RAND_1189[7:0];
  _RAND_1190 = {1{`RANDOM}};
  frameBuffer_9_22 = _RAND_1190[7:0];
  _RAND_1191 = {1{`RANDOM}};
  frameBuffer_9_23 = _RAND_1191[7:0];
  _RAND_1192 = {1{`RANDOM}};
  frameBuffer_9_24 = _RAND_1192[7:0];
  _RAND_1193 = {1{`RANDOM}};
  frameBuffer_9_25 = _RAND_1193[7:0];
  _RAND_1194 = {1{`RANDOM}};
  frameBuffer_9_26 = _RAND_1194[7:0];
  _RAND_1195 = {1{`RANDOM}};
  frameBuffer_9_27 = _RAND_1195[7:0];
  _RAND_1196 = {1{`RANDOM}};
  frameBuffer_9_28 = _RAND_1196[7:0];
  _RAND_1197 = {1{`RANDOM}};
  frameBuffer_9_29 = _RAND_1197[7:0];
  _RAND_1198 = {1{`RANDOM}};
  frameBuffer_9_30 = _RAND_1198[7:0];
  _RAND_1199 = {1{`RANDOM}};
  frameBuffer_9_31 = _RAND_1199[7:0];
  _RAND_1200 = {1{`RANDOM}};
  frameBuffer_9_32 = _RAND_1200[7:0];
  _RAND_1201 = {1{`RANDOM}};
  frameBuffer_9_33 = _RAND_1201[7:0];
  _RAND_1202 = {1{`RANDOM}};
  frameBuffer_9_34 = _RAND_1202[7:0];
  _RAND_1203 = {1{`RANDOM}};
  frameBuffer_9_35 = _RAND_1203[7:0];
  _RAND_1204 = {1{`RANDOM}};
  frameBuffer_9_36 = _RAND_1204[7:0];
  _RAND_1205 = {1{`RANDOM}};
  frameBuffer_9_37 = _RAND_1205[7:0];
  _RAND_1206 = {1{`RANDOM}};
  frameBuffer_9_38 = _RAND_1206[7:0];
  _RAND_1207 = {1{`RANDOM}};
  frameBuffer_9_39 = _RAND_1207[7:0];
  _RAND_1208 = {1{`RANDOM}};
  frameBuffer_9_40 = _RAND_1208[7:0];
  _RAND_1209 = {1{`RANDOM}};
  frameBuffer_9_41 = _RAND_1209[7:0];
  _RAND_1210 = {1{`RANDOM}};
  frameBuffer_9_42 = _RAND_1210[7:0];
  _RAND_1211 = {1{`RANDOM}};
  frameBuffer_9_43 = _RAND_1211[7:0];
  _RAND_1212 = {1{`RANDOM}};
  frameBuffer_9_44 = _RAND_1212[7:0];
  _RAND_1213 = {1{`RANDOM}};
  frameBuffer_9_45 = _RAND_1213[7:0];
  _RAND_1214 = {1{`RANDOM}};
  frameBuffer_9_46 = _RAND_1214[7:0];
  _RAND_1215 = {1{`RANDOM}};
  frameBuffer_9_47 = _RAND_1215[7:0];
  _RAND_1216 = {1{`RANDOM}};
  frameBuffer_9_48 = _RAND_1216[7:0];
  _RAND_1217 = {1{`RANDOM}};
  frameBuffer_9_49 = _RAND_1217[7:0];
  _RAND_1218 = {1{`RANDOM}};
  frameBuffer_9_50 = _RAND_1218[7:0];
  _RAND_1219 = {1{`RANDOM}};
  frameBuffer_9_51 = _RAND_1219[7:0];
  _RAND_1220 = {1{`RANDOM}};
  frameBuffer_9_52 = _RAND_1220[7:0];
  _RAND_1221 = {1{`RANDOM}};
  frameBuffer_9_53 = _RAND_1221[7:0];
  _RAND_1222 = {1{`RANDOM}};
  frameBuffer_9_54 = _RAND_1222[7:0];
  _RAND_1223 = {1{`RANDOM}};
  frameBuffer_9_55 = _RAND_1223[7:0];
  _RAND_1224 = {1{`RANDOM}};
  frameBuffer_9_56 = _RAND_1224[7:0];
  _RAND_1225 = {1{`RANDOM}};
  frameBuffer_9_57 = _RAND_1225[7:0];
  _RAND_1226 = {1{`RANDOM}};
  frameBuffer_9_58 = _RAND_1226[7:0];
  _RAND_1227 = {1{`RANDOM}};
  frameBuffer_9_59 = _RAND_1227[7:0];
  _RAND_1228 = {1{`RANDOM}};
  frameBuffer_9_60 = _RAND_1228[7:0];
  _RAND_1229 = {1{`RANDOM}};
  frameBuffer_9_61 = _RAND_1229[7:0];
  _RAND_1230 = {1{`RANDOM}};
  frameBuffer_9_62 = _RAND_1230[7:0];
  _RAND_1231 = {1{`RANDOM}};
  frameBuffer_9_63 = _RAND_1231[7:0];
  _RAND_1232 = {1{`RANDOM}};
  frameBuffer_9_64 = _RAND_1232[7:0];
  _RAND_1233 = {1{`RANDOM}};
  frameBuffer_9_65 = _RAND_1233[7:0];
  _RAND_1234 = {1{`RANDOM}};
  frameBuffer_9_66 = _RAND_1234[7:0];
  _RAND_1235 = {1{`RANDOM}};
  frameBuffer_9_67 = _RAND_1235[7:0];
  _RAND_1236 = {1{`RANDOM}};
  frameBuffer_9_68 = _RAND_1236[7:0];
  _RAND_1237 = {1{`RANDOM}};
  frameBuffer_9_69 = _RAND_1237[7:0];
  _RAND_1238 = {1{`RANDOM}};
  frameBuffer_9_70 = _RAND_1238[7:0];
  _RAND_1239 = {1{`RANDOM}};
  frameBuffer_9_71 = _RAND_1239[7:0];
  _RAND_1240 = {1{`RANDOM}};
  frameBuffer_9_72 = _RAND_1240[7:0];
  _RAND_1241 = {1{`RANDOM}};
  frameBuffer_9_73 = _RAND_1241[7:0];
  _RAND_1242 = {1{`RANDOM}};
  frameBuffer_9_74 = _RAND_1242[7:0];
  _RAND_1243 = {1{`RANDOM}};
  frameBuffer_9_75 = _RAND_1243[7:0];
  _RAND_1244 = {1{`RANDOM}};
  frameBuffer_9_76 = _RAND_1244[7:0];
  _RAND_1245 = {1{`RANDOM}};
  frameBuffer_9_77 = _RAND_1245[7:0];
  _RAND_1246 = {1{`RANDOM}};
  frameBuffer_9_78 = _RAND_1246[7:0];
  _RAND_1247 = {1{`RANDOM}};
  frameBuffer_9_79 = _RAND_1247[7:0];
  _RAND_1248 = {1{`RANDOM}};
  frameBuffer_9_80 = _RAND_1248[7:0];
  _RAND_1249 = {1{`RANDOM}};
  frameBuffer_9_81 = _RAND_1249[7:0];
  _RAND_1250 = {1{`RANDOM}};
  frameBuffer_9_82 = _RAND_1250[7:0];
  _RAND_1251 = {1{`RANDOM}};
  frameBuffer_9_83 = _RAND_1251[7:0];
  _RAND_1252 = {1{`RANDOM}};
  frameBuffer_9_84 = _RAND_1252[7:0];
  _RAND_1253 = {1{`RANDOM}};
  frameBuffer_9_85 = _RAND_1253[7:0];
  _RAND_1254 = {1{`RANDOM}};
  frameBuffer_9_86 = _RAND_1254[7:0];
  _RAND_1255 = {1{`RANDOM}};
  frameBuffer_9_87 = _RAND_1255[7:0];
  _RAND_1256 = {1{`RANDOM}};
  frameBuffer_9_88 = _RAND_1256[7:0];
  _RAND_1257 = {1{`RANDOM}};
  frameBuffer_9_89 = _RAND_1257[7:0];
  _RAND_1258 = {1{`RANDOM}};
  frameBuffer_9_90 = _RAND_1258[7:0];
  _RAND_1259 = {1{`RANDOM}};
  frameBuffer_9_91 = _RAND_1259[7:0];
  _RAND_1260 = {1{`RANDOM}};
  frameBuffer_9_92 = _RAND_1260[7:0];
  _RAND_1261 = {1{`RANDOM}};
  frameBuffer_9_93 = _RAND_1261[7:0];
  _RAND_1262 = {1{`RANDOM}};
  frameBuffer_9_94 = _RAND_1262[7:0];
  _RAND_1263 = {1{`RANDOM}};
  frameBuffer_9_95 = _RAND_1263[7:0];
  _RAND_1264 = {1{`RANDOM}};
  frameBuffer_9_96 = _RAND_1264[7:0];
  _RAND_1265 = {1{`RANDOM}};
  frameBuffer_9_97 = _RAND_1265[7:0];
  _RAND_1266 = {1{`RANDOM}};
  frameBuffer_9_98 = _RAND_1266[7:0];
  _RAND_1267 = {1{`RANDOM}};
  frameBuffer_9_99 = _RAND_1267[7:0];
  _RAND_1268 = {1{`RANDOM}};
  frameBuffer_9_100 = _RAND_1268[7:0];
  _RAND_1269 = {1{`RANDOM}};
  frameBuffer_9_101 = _RAND_1269[7:0];
  _RAND_1270 = {1{`RANDOM}};
  frameBuffer_9_102 = _RAND_1270[7:0];
  _RAND_1271 = {1{`RANDOM}};
  frameBuffer_9_103 = _RAND_1271[7:0];
  _RAND_1272 = {1{`RANDOM}};
  frameBuffer_9_104 = _RAND_1272[7:0];
  _RAND_1273 = {1{`RANDOM}};
  frameBuffer_9_105 = _RAND_1273[7:0];
  _RAND_1274 = {1{`RANDOM}};
  frameBuffer_9_106 = _RAND_1274[7:0];
  _RAND_1275 = {1{`RANDOM}};
  frameBuffer_9_107 = _RAND_1275[7:0];
  _RAND_1276 = {1{`RANDOM}};
  frameBuffer_9_108 = _RAND_1276[7:0];
  _RAND_1277 = {1{`RANDOM}};
  frameBuffer_9_109 = _RAND_1277[7:0];
  _RAND_1278 = {1{`RANDOM}};
  frameBuffer_9_110 = _RAND_1278[7:0];
  _RAND_1279 = {1{`RANDOM}};
  frameBuffer_9_111 = _RAND_1279[7:0];
  _RAND_1280 = {1{`RANDOM}};
  frameBuffer_9_112 = _RAND_1280[7:0];
  _RAND_1281 = {1{`RANDOM}};
  frameBuffer_9_113 = _RAND_1281[7:0];
  _RAND_1282 = {1{`RANDOM}};
  frameBuffer_9_114 = _RAND_1282[7:0];
  _RAND_1283 = {1{`RANDOM}};
  frameBuffer_9_115 = _RAND_1283[7:0];
  _RAND_1284 = {1{`RANDOM}};
  frameBuffer_9_116 = _RAND_1284[7:0];
  _RAND_1285 = {1{`RANDOM}};
  frameBuffer_9_117 = _RAND_1285[7:0];
  _RAND_1286 = {1{`RANDOM}};
  frameBuffer_9_118 = _RAND_1286[7:0];
  _RAND_1287 = {1{`RANDOM}};
  frameBuffer_9_119 = _RAND_1287[7:0];
  _RAND_1288 = {1{`RANDOM}};
  frameBuffer_9_120 = _RAND_1288[7:0];
  _RAND_1289 = {1{`RANDOM}};
  frameBuffer_9_121 = _RAND_1289[7:0];
  _RAND_1290 = {1{`RANDOM}};
  frameBuffer_9_122 = _RAND_1290[7:0];
  _RAND_1291 = {1{`RANDOM}};
  frameBuffer_9_123 = _RAND_1291[7:0];
  _RAND_1292 = {1{`RANDOM}};
  frameBuffer_9_124 = _RAND_1292[7:0];
  _RAND_1293 = {1{`RANDOM}};
  frameBuffer_9_125 = _RAND_1293[7:0];
  _RAND_1294 = {1{`RANDOM}};
  frameBuffer_9_126 = _RAND_1294[7:0];
  _RAND_1295 = {1{`RANDOM}};
  frameBuffer_9_127 = _RAND_1295[7:0];
  _RAND_1296 = {1{`RANDOM}};
  frameBuffer_10_0 = _RAND_1296[7:0];
  _RAND_1297 = {1{`RANDOM}};
  frameBuffer_10_1 = _RAND_1297[7:0];
  _RAND_1298 = {1{`RANDOM}};
  frameBuffer_10_2 = _RAND_1298[7:0];
  _RAND_1299 = {1{`RANDOM}};
  frameBuffer_10_3 = _RAND_1299[7:0];
  _RAND_1300 = {1{`RANDOM}};
  frameBuffer_10_4 = _RAND_1300[7:0];
  _RAND_1301 = {1{`RANDOM}};
  frameBuffer_10_5 = _RAND_1301[7:0];
  _RAND_1302 = {1{`RANDOM}};
  frameBuffer_10_6 = _RAND_1302[7:0];
  _RAND_1303 = {1{`RANDOM}};
  frameBuffer_10_7 = _RAND_1303[7:0];
  _RAND_1304 = {1{`RANDOM}};
  frameBuffer_10_8 = _RAND_1304[7:0];
  _RAND_1305 = {1{`RANDOM}};
  frameBuffer_10_9 = _RAND_1305[7:0];
  _RAND_1306 = {1{`RANDOM}};
  frameBuffer_10_10 = _RAND_1306[7:0];
  _RAND_1307 = {1{`RANDOM}};
  frameBuffer_10_11 = _RAND_1307[7:0];
  _RAND_1308 = {1{`RANDOM}};
  frameBuffer_10_12 = _RAND_1308[7:0];
  _RAND_1309 = {1{`RANDOM}};
  frameBuffer_10_13 = _RAND_1309[7:0];
  _RAND_1310 = {1{`RANDOM}};
  frameBuffer_10_14 = _RAND_1310[7:0];
  _RAND_1311 = {1{`RANDOM}};
  frameBuffer_10_15 = _RAND_1311[7:0];
  _RAND_1312 = {1{`RANDOM}};
  frameBuffer_10_16 = _RAND_1312[7:0];
  _RAND_1313 = {1{`RANDOM}};
  frameBuffer_10_17 = _RAND_1313[7:0];
  _RAND_1314 = {1{`RANDOM}};
  frameBuffer_10_18 = _RAND_1314[7:0];
  _RAND_1315 = {1{`RANDOM}};
  frameBuffer_10_19 = _RAND_1315[7:0];
  _RAND_1316 = {1{`RANDOM}};
  frameBuffer_10_20 = _RAND_1316[7:0];
  _RAND_1317 = {1{`RANDOM}};
  frameBuffer_10_21 = _RAND_1317[7:0];
  _RAND_1318 = {1{`RANDOM}};
  frameBuffer_10_22 = _RAND_1318[7:0];
  _RAND_1319 = {1{`RANDOM}};
  frameBuffer_10_23 = _RAND_1319[7:0];
  _RAND_1320 = {1{`RANDOM}};
  frameBuffer_10_24 = _RAND_1320[7:0];
  _RAND_1321 = {1{`RANDOM}};
  frameBuffer_10_25 = _RAND_1321[7:0];
  _RAND_1322 = {1{`RANDOM}};
  frameBuffer_10_26 = _RAND_1322[7:0];
  _RAND_1323 = {1{`RANDOM}};
  frameBuffer_10_27 = _RAND_1323[7:0];
  _RAND_1324 = {1{`RANDOM}};
  frameBuffer_10_28 = _RAND_1324[7:0];
  _RAND_1325 = {1{`RANDOM}};
  frameBuffer_10_29 = _RAND_1325[7:0];
  _RAND_1326 = {1{`RANDOM}};
  frameBuffer_10_30 = _RAND_1326[7:0];
  _RAND_1327 = {1{`RANDOM}};
  frameBuffer_10_31 = _RAND_1327[7:0];
  _RAND_1328 = {1{`RANDOM}};
  frameBuffer_10_32 = _RAND_1328[7:0];
  _RAND_1329 = {1{`RANDOM}};
  frameBuffer_10_33 = _RAND_1329[7:0];
  _RAND_1330 = {1{`RANDOM}};
  frameBuffer_10_34 = _RAND_1330[7:0];
  _RAND_1331 = {1{`RANDOM}};
  frameBuffer_10_35 = _RAND_1331[7:0];
  _RAND_1332 = {1{`RANDOM}};
  frameBuffer_10_36 = _RAND_1332[7:0];
  _RAND_1333 = {1{`RANDOM}};
  frameBuffer_10_37 = _RAND_1333[7:0];
  _RAND_1334 = {1{`RANDOM}};
  frameBuffer_10_38 = _RAND_1334[7:0];
  _RAND_1335 = {1{`RANDOM}};
  frameBuffer_10_39 = _RAND_1335[7:0];
  _RAND_1336 = {1{`RANDOM}};
  frameBuffer_10_40 = _RAND_1336[7:0];
  _RAND_1337 = {1{`RANDOM}};
  frameBuffer_10_41 = _RAND_1337[7:0];
  _RAND_1338 = {1{`RANDOM}};
  frameBuffer_10_42 = _RAND_1338[7:0];
  _RAND_1339 = {1{`RANDOM}};
  frameBuffer_10_43 = _RAND_1339[7:0];
  _RAND_1340 = {1{`RANDOM}};
  frameBuffer_10_44 = _RAND_1340[7:0];
  _RAND_1341 = {1{`RANDOM}};
  frameBuffer_10_45 = _RAND_1341[7:0];
  _RAND_1342 = {1{`RANDOM}};
  frameBuffer_10_46 = _RAND_1342[7:0];
  _RAND_1343 = {1{`RANDOM}};
  frameBuffer_10_47 = _RAND_1343[7:0];
  _RAND_1344 = {1{`RANDOM}};
  frameBuffer_10_48 = _RAND_1344[7:0];
  _RAND_1345 = {1{`RANDOM}};
  frameBuffer_10_49 = _RAND_1345[7:0];
  _RAND_1346 = {1{`RANDOM}};
  frameBuffer_10_50 = _RAND_1346[7:0];
  _RAND_1347 = {1{`RANDOM}};
  frameBuffer_10_51 = _RAND_1347[7:0];
  _RAND_1348 = {1{`RANDOM}};
  frameBuffer_10_52 = _RAND_1348[7:0];
  _RAND_1349 = {1{`RANDOM}};
  frameBuffer_10_53 = _RAND_1349[7:0];
  _RAND_1350 = {1{`RANDOM}};
  frameBuffer_10_54 = _RAND_1350[7:0];
  _RAND_1351 = {1{`RANDOM}};
  frameBuffer_10_55 = _RAND_1351[7:0];
  _RAND_1352 = {1{`RANDOM}};
  frameBuffer_10_56 = _RAND_1352[7:0];
  _RAND_1353 = {1{`RANDOM}};
  frameBuffer_10_57 = _RAND_1353[7:0];
  _RAND_1354 = {1{`RANDOM}};
  frameBuffer_10_58 = _RAND_1354[7:0];
  _RAND_1355 = {1{`RANDOM}};
  frameBuffer_10_59 = _RAND_1355[7:0];
  _RAND_1356 = {1{`RANDOM}};
  frameBuffer_10_60 = _RAND_1356[7:0];
  _RAND_1357 = {1{`RANDOM}};
  frameBuffer_10_61 = _RAND_1357[7:0];
  _RAND_1358 = {1{`RANDOM}};
  frameBuffer_10_62 = _RAND_1358[7:0];
  _RAND_1359 = {1{`RANDOM}};
  frameBuffer_10_63 = _RAND_1359[7:0];
  _RAND_1360 = {1{`RANDOM}};
  frameBuffer_10_64 = _RAND_1360[7:0];
  _RAND_1361 = {1{`RANDOM}};
  frameBuffer_10_65 = _RAND_1361[7:0];
  _RAND_1362 = {1{`RANDOM}};
  frameBuffer_10_66 = _RAND_1362[7:0];
  _RAND_1363 = {1{`RANDOM}};
  frameBuffer_10_67 = _RAND_1363[7:0];
  _RAND_1364 = {1{`RANDOM}};
  frameBuffer_10_68 = _RAND_1364[7:0];
  _RAND_1365 = {1{`RANDOM}};
  frameBuffer_10_69 = _RAND_1365[7:0];
  _RAND_1366 = {1{`RANDOM}};
  frameBuffer_10_70 = _RAND_1366[7:0];
  _RAND_1367 = {1{`RANDOM}};
  frameBuffer_10_71 = _RAND_1367[7:0];
  _RAND_1368 = {1{`RANDOM}};
  frameBuffer_10_72 = _RAND_1368[7:0];
  _RAND_1369 = {1{`RANDOM}};
  frameBuffer_10_73 = _RAND_1369[7:0];
  _RAND_1370 = {1{`RANDOM}};
  frameBuffer_10_74 = _RAND_1370[7:0];
  _RAND_1371 = {1{`RANDOM}};
  frameBuffer_10_75 = _RAND_1371[7:0];
  _RAND_1372 = {1{`RANDOM}};
  frameBuffer_10_76 = _RAND_1372[7:0];
  _RAND_1373 = {1{`RANDOM}};
  frameBuffer_10_77 = _RAND_1373[7:0];
  _RAND_1374 = {1{`RANDOM}};
  frameBuffer_10_78 = _RAND_1374[7:0];
  _RAND_1375 = {1{`RANDOM}};
  frameBuffer_10_79 = _RAND_1375[7:0];
  _RAND_1376 = {1{`RANDOM}};
  frameBuffer_10_80 = _RAND_1376[7:0];
  _RAND_1377 = {1{`RANDOM}};
  frameBuffer_10_81 = _RAND_1377[7:0];
  _RAND_1378 = {1{`RANDOM}};
  frameBuffer_10_82 = _RAND_1378[7:0];
  _RAND_1379 = {1{`RANDOM}};
  frameBuffer_10_83 = _RAND_1379[7:0];
  _RAND_1380 = {1{`RANDOM}};
  frameBuffer_10_84 = _RAND_1380[7:0];
  _RAND_1381 = {1{`RANDOM}};
  frameBuffer_10_85 = _RAND_1381[7:0];
  _RAND_1382 = {1{`RANDOM}};
  frameBuffer_10_86 = _RAND_1382[7:0];
  _RAND_1383 = {1{`RANDOM}};
  frameBuffer_10_87 = _RAND_1383[7:0];
  _RAND_1384 = {1{`RANDOM}};
  frameBuffer_10_88 = _RAND_1384[7:0];
  _RAND_1385 = {1{`RANDOM}};
  frameBuffer_10_89 = _RAND_1385[7:0];
  _RAND_1386 = {1{`RANDOM}};
  frameBuffer_10_90 = _RAND_1386[7:0];
  _RAND_1387 = {1{`RANDOM}};
  frameBuffer_10_91 = _RAND_1387[7:0];
  _RAND_1388 = {1{`RANDOM}};
  frameBuffer_10_92 = _RAND_1388[7:0];
  _RAND_1389 = {1{`RANDOM}};
  frameBuffer_10_93 = _RAND_1389[7:0];
  _RAND_1390 = {1{`RANDOM}};
  frameBuffer_10_94 = _RAND_1390[7:0];
  _RAND_1391 = {1{`RANDOM}};
  frameBuffer_10_95 = _RAND_1391[7:0];
  _RAND_1392 = {1{`RANDOM}};
  frameBuffer_10_96 = _RAND_1392[7:0];
  _RAND_1393 = {1{`RANDOM}};
  frameBuffer_10_97 = _RAND_1393[7:0];
  _RAND_1394 = {1{`RANDOM}};
  frameBuffer_10_98 = _RAND_1394[7:0];
  _RAND_1395 = {1{`RANDOM}};
  frameBuffer_10_99 = _RAND_1395[7:0];
  _RAND_1396 = {1{`RANDOM}};
  frameBuffer_10_100 = _RAND_1396[7:0];
  _RAND_1397 = {1{`RANDOM}};
  frameBuffer_10_101 = _RAND_1397[7:0];
  _RAND_1398 = {1{`RANDOM}};
  frameBuffer_10_102 = _RAND_1398[7:0];
  _RAND_1399 = {1{`RANDOM}};
  frameBuffer_10_103 = _RAND_1399[7:0];
  _RAND_1400 = {1{`RANDOM}};
  frameBuffer_10_104 = _RAND_1400[7:0];
  _RAND_1401 = {1{`RANDOM}};
  frameBuffer_10_105 = _RAND_1401[7:0];
  _RAND_1402 = {1{`RANDOM}};
  frameBuffer_10_106 = _RAND_1402[7:0];
  _RAND_1403 = {1{`RANDOM}};
  frameBuffer_10_107 = _RAND_1403[7:0];
  _RAND_1404 = {1{`RANDOM}};
  frameBuffer_10_108 = _RAND_1404[7:0];
  _RAND_1405 = {1{`RANDOM}};
  frameBuffer_10_109 = _RAND_1405[7:0];
  _RAND_1406 = {1{`RANDOM}};
  frameBuffer_10_110 = _RAND_1406[7:0];
  _RAND_1407 = {1{`RANDOM}};
  frameBuffer_10_111 = _RAND_1407[7:0];
  _RAND_1408 = {1{`RANDOM}};
  frameBuffer_10_112 = _RAND_1408[7:0];
  _RAND_1409 = {1{`RANDOM}};
  frameBuffer_10_113 = _RAND_1409[7:0];
  _RAND_1410 = {1{`RANDOM}};
  frameBuffer_10_114 = _RAND_1410[7:0];
  _RAND_1411 = {1{`RANDOM}};
  frameBuffer_10_115 = _RAND_1411[7:0];
  _RAND_1412 = {1{`RANDOM}};
  frameBuffer_10_116 = _RAND_1412[7:0];
  _RAND_1413 = {1{`RANDOM}};
  frameBuffer_10_117 = _RAND_1413[7:0];
  _RAND_1414 = {1{`RANDOM}};
  frameBuffer_10_118 = _RAND_1414[7:0];
  _RAND_1415 = {1{`RANDOM}};
  frameBuffer_10_119 = _RAND_1415[7:0];
  _RAND_1416 = {1{`RANDOM}};
  frameBuffer_10_120 = _RAND_1416[7:0];
  _RAND_1417 = {1{`RANDOM}};
  frameBuffer_10_121 = _RAND_1417[7:0];
  _RAND_1418 = {1{`RANDOM}};
  frameBuffer_10_122 = _RAND_1418[7:0];
  _RAND_1419 = {1{`RANDOM}};
  frameBuffer_10_123 = _RAND_1419[7:0];
  _RAND_1420 = {1{`RANDOM}};
  frameBuffer_10_124 = _RAND_1420[7:0];
  _RAND_1421 = {1{`RANDOM}};
  frameBuffer_10_125 = _RAND_1421[7:0];
  _RAND_1422 = {1{`RANDOM}};
  frameBuffer_10_126 = _RAND_1422[7:0];
  _RAND_1423 = {1{`RANDOM}};
  frameBuffer_10_127 = _RAND_1423[7:0];
  _RAND_1424 = {1{`RANDOM}};
  frameBuffer_11_0 = _RAND_1424[7:0];
  _RAND_1425 = {1{`RANDOM}};
  frameBuffer_11_1 = _RAND_1425[7:0];
  _RAND_1426 = {1{`RANDOM}};
  frameBuffer_11_2 = _RAND_1426[7:0];
  _RAND_1427 = {1{`RANDOM}};
  frameBuffer_11_3 = _RAND_1427[7:0];
  _RAND_1428 = {1{`RANDOM}};
  frameBuffer_11_4 = _RAND_1428[7:0];
  _RAND_1429 = {1{`RANDOM}};
  frameBuffer_11_5 = _RAND_1429[7:0];
  _RAND_1430 = {1{`RANDOM}};
  frameBuffer_11_6 = _RAND_1430[7:0];
  _RAND_1431 = {1{`RANDOM}};
  frameBuffer_11_7 = _RAND_1431[7:0];
  _RAND_1432 = {1{`RANDOM}};
  frameBuffer_11_8 = _RAND_1432[7:0];
  _RAND_1433 = {1{`RANDOM}};
  frameBuffer_11_9 = _RAND_1433[7:0];
  _RAND_1434 = {1{`RANDOM}};
  frameBuffer_11_10 = _RAND_1434[7:0];
  _RAND_1435 = {1{`RANDOM}};
  frameBuffer_11_11 = _RAND_1435[7:0];
  _RAND_1436 = {1{`RANDOM}};
  frameBuffer_11_12 = _RAND_1436[7:0];
  _RAND_1437 = {1{`RANDOM}};
  frameBuffer_11_13 = _RAND_1437[7:0];
  _RAND_1438 = {1{`RANDOM}};
  frameBuffer_11_14 = _RAND_1438[7:0];
  _RAND_1439 = {1{`RANDOM}};
  frameBuffer_11_15 = _RAND_1439[7:0];
  _RAND_1440 = {1{`RANDOM}};
  frameBuffer_11_16 = _RAND_1440[7:0];
  _RAND_1441 = {1{`RANDOM}};
  frameBuffer_11_17 = _RAND_1441[7:0];
  _RAND_1442 = {1{`RANDOM}};
  frameBuffer_11_18 = _RAND_1442[7:0];
  _RAND_1443 = {1{`RANDOM}};
  frameBuffer_11_19 = _RAND_1443[7:0];
  _RAND_1444 = {1{`RANDOM}};
  frameBuffer_11_20 = _RAND_1444[7:0];
  _RAND_1445 = {1{`RANDOM}};
  frameBuffer_11_21 = _RAND_1445[7:0];
  _RAND_1446 = {1{`RANDOM}};
  frameBuffer_11_22 = _RAND_1446[7:0];
  _RAND_1447 = {1{`RANDOM}};
  frameBuffer_11_23 = _RAND_1447[7:0];
  _RAND_1448 = {1{`RANDOM}};
  frameBuffer_11_24 = _RAND_1448[7:0];
  _RAND_1449 = {1{`RANDOM}};
  frameBuffer_11_25 = _RAND_1449[7:0];
  _RAND_1450 = {1{`RANDOM}};
  frameBuffer_11_26 = _RAND_1450[7:0];
  _RAND_1451 = {1{`RANDOM}};
  frameBuffer_11_27 = _RAND_1451[7:0];
  _RAND_1452 = {1{`RANDOM}};
  frameBuffer_11_28 = _RAND_1452[7:0];
  _RAND_1453 = {1{`RANDOM}};
  frameBuffer_11_29 = _RAND_1453[7:0];
  _RAND_1454 = {1{`RANDOM}};
  frameBuffer_11_30 = _RAND_1454[7:0];
  _RAND_1455 = {1{`RANDOM}};
  frameBuffer_11_31 = _RAND_1455[7:0];
  _RAND_1456 = {1{`RANDOM}};
  frameBuffer_11_32 = _RAND_1456[7:0];
  _RAND_1457 = {1{`RANDOM}};
  frameBuffer_11_33 = _RAND_1457[7:0];
  _RAND_1458 = {1{`RANDOM}};
  frameBuffer_11_34 = _RAND_1458[7:0];
  _RAND_1459 = {1{`RANDOM}};
  frameBuffer_11_35 = _RAND_1459[7:0];
  _RAND_1460 = {1{`RANDOM}};
  frameBuffer_11_36 = _RAND_1460[7:0];
  _RAND_1461 = {1{`RANDOM}};
  frameBuffer_11_37 = _RAND_1461[7:0];
  _RAND_1462 = {1{`RANDOM}};
  frameBuffer_11_38 = _RAND_1462[7:0];
  _RAND_1463 = {1{`RANDOM}};
  frameBuffer_11_39 = _RAND_1463[7:0];
  _RAND_1464 = {1{`RANDOM}};
  frameBuffer_11_40 = _RAND_1464[7:0];
  _RAND_1465 = {1{`RANDOM}};
  frameBuffer_11_41 = _RAND_1465[7:0];
  _RAND_1466 = {1{`RANDOM}};
  frameBuffer_11_42 = _RAND_1466[7:0];
  _RAND_1467 = {1{`RANDOM}};
  frameBuffer_11_43 = _RAND_1467[7:0];
  _RAND_1468 = {1{`RANDOM}};
  frameBuffer_11_44 = _RAND_1468[7:0];
  _RAND_1469 = {1{`RANDOM}};
  frameBuffer_11_45 = _RAND_1469[7:0];
  _RAND_1470 = {1{`RANDOM}};
  frameBuffer_11_46 = _RAND_1470[7:0];
  _RAND_1471 = {1{`RANDOM}};
  frameBuffer_11_47 = _RAND_1471[7:0];
  _RAND_1472 = {1{`RANDOM}};
  frameBuffer_11_48 = _RAND_1472[7:0];
  _RAND_1473 = {1{`RANDOM}};
  frameBuffer_11_49 = _RAND_1473[7:0];
  _RAND_1474 = {1{`RANDOM}};
  frameBuffer_11_50 = _RAND_1474[7:0];
  _RAND_1475 = {1{`RANDOM}};
  frameBuffer_11_51 = _RAND_1475[7:0];
  _RAND_1476 = {1{`RANDOM}};
  frameBuffer_11_52 = _RAND_1476[7:0];
  _RAND_1477 = {1{`RANDOM}};
  frameBuffer_11_53 = _RAND_1477[7:0];
  _RAND_1478 = {1{`RANDOM}};
  frameBuffer_11_54 = _RAND_1478[7:0];
  _RAND_1479 = {1{`RANDOM}};
  frameBuffer_11_55 = _RAND_1479[7:0];
  _RAND_1480 = {1{`RANDOM}};
  frameBuffer_11_56 = _RAND_1480[7:0];
  _RAND_1481 = {1{`RANDOM}};
  frameBuffer_11_57 = _RAND_1481[7:0];
  _RAND_1482 = {1{`RANDOM}};
  frameBuffer_11_58 = _RAND_1482[7:0];
  _RAND_1483 = {1{`RANDOM}};
  frameBuffer_11_59 = _RAND_1483[7:0];
  _RAND_1484 = {1{`RANDOM}};
  frameBuffer_11_60 = _RAND_1484[7:0];
  _RAND_1485 = {1{`RANDOM}};
  frameBuffer_11_61 = _RAND_1485[7:0];
  _RAND_1486 = {1{`RANDOM}};
  frameBuffer_11_62 = _RAND_1486[7:0];
  _RAND_1487 = {1{`RANDOM}};
  frameBuffer_11_63 = _RAND_1487[7:0];
  _RAND_1488 = {1{`RANDOM}};
  frameBuffer_11_64 = _RAND_1488[7:0];
  _RAND_1489 = {1{`RANDOM}};
  frameBuffer_11_65 = _RAND_1489[7:0];
  _RAND_1490 = {1{`RANDOM}};
  frameBuffer_11_66 = _RAND_1490[7:0];
  _RAND_1491 = {1{`RANDOM}};
  frameBuffer_11_67 = _RAND_1491[7:0];
  _RAND_1492 = {1{`RANDOM}};
  frameBuffer_11_68 = _RAND_1492[7:0];
  _RAND_1493 = {1{`RANDOM}};
  frameBuffer_11_69 = _RAND_1493[7:0];
  _RAND_1494 = {1{`RANDOM}};
  frameBuffer_11_70 = _RAND_1494[7:0];
  _RAND_1495 = {1{`RANDOM}};
  frameBuffer_11_71 = _RAND_1495[7:0];
  _RAND_1496 = {1{`RANDOM}};
  frameBuffer_11_72 = _RAND_1496[7:0];
  _RAND_1497 = {1{`RANDOM}};
  frameBuffer_11_73 = _RAND_1497[7:0];
  _RAND_1498 = {1{`RANDOM}};
  frameBuffer_11_74 = _RAND_1498[7:0];
  _RAND_1499 = {1{`RANDOM}};
  frameBuffer_11_75 = _RAND_1499[7:0];
  _RAND_1500 = {1{`RANDOM}};
  frameBuffer_11_76 = _RAND_1500[7:0];
  _RAND_1501 = {1{`RANDOM}};
  frameBuffer_11_77 = _RAND_1501[7:0];
  _RAND_1502 = {1{`RANDOM}};
  frameBuffer_11_78 = _RAND_1502[7:0];
  _RAND_1503 = {1{`RANDOM}};
  frameBuffer_11_79 = _RAND_1503[7:0];
  _RAND_1504 = {1{`RANDOM}};
  frameBuffer_11_80 = _RAND_1504[7:0];
  _RAND_1505 = {1{`RANDOM}};
  frameBuffer_11_81 = _RAND_1505[7:0];
  _RAND_1506 = {1{`RANDOM}};
  frameBuffer_11_82 = _RAND_1506[7:0];
  _RAND_1507 = {1{`RANDOM}};
  frameBuffer_11_83 = _RAND_1507[7:0];
  _RAND_1508 = {1{`RANDOM}};
  frameBuffer_11_84 = _RAND_1508[7:0];
  _RAND_1509 = {1{`RANDOM}};
  frameBuffer_11_85 = _RAND_1509[7:0];
  _RAND_1510 = {1{`RANDOM}};
  frameBuffer_11_86 = _RAND_1510[7:0];
  _RAND_1511 = {1{`RANDOM}};
  frameBuffer_11_87 = _RAND_1511[7:0];
  _RAND_1512 = {1{`RANDOM}};
  frameBuffer_11_88 = _RAND_1512[7:0];
  _RAND_1513 = {1{`RANDOM}};
  frameBuffer_11_89 = _RAND_1513[7:0];
  _RAND_1514 = {1{`RANDOM}};
  frameBuffer_11_90 = _RAND_1514[7:0];
  _RAND_1515 = {1{`RANDOM}};
  frameBuffer_11_91 = _RAND_1515[7:0];
  _RAND_1516 = {1{`RANDOM}};
  frameBuffer_11_92 = _RAND_1516[7:0];
  _RAND_1517 = {1{`RANDOM}};
  frameBuffer_11_93 = _RAND_1517[7:0];
  _RAND_1518 = {1{`RANDOM}};
  frameBuffer_11_94 = _RAND_1518[7:0];
  _RAND_1519 = {1{`RANDOM}};
  frameBuffer_11_95 = _RAND_1519[7:0];
  _RAND_1520 = {1{`RANDOM}};
  frameBuffer_11_96 = _RAND_1520[7:0];
  _RAND_1521 = {1{`RANDOM}};
  frameBuffer_11_97 = _RAND_1521[7:0];
  _RAND_1522 = {1{`RANDOM}};
  frameBuffer_11_98 = _RAND_1522[7:0];
  _RAND_1523 = {1{`RANDOM}};
  frameBuffer_11_99 = _RAND_1523[7:0];
  _RAND_1524 = {1{`RANDOM}};
  frameBuffer_11_100 = _RAND_1524[7:0];
  _RAND_1525 = {1{`RANDOM}};
  frameBuffer_11_101 = _RAND_1525[7:0];
  _RAND_1526 = {1{`RANDOM}};
  frameBuffer_11_102 = _RAND_1526[7:0];
  _RAND_1527 = {1{`RANDOM}};
  frameBuffer_11_103 = _RAND_1527[7:0];
  _RAND_1528 = {1{`RANDOM}};
  frameBuffer_11_104 = _RAND_1528[7:0];
  _RAND_1529 = {1{`RANDOM}};
  frameBuffer_11_105 = _RAND_1529[7:0];
  _RAND_1530 = {1{`RANDOM}};
  frameBuffer_11_106 = _RAND_1530[7:0];
  _RAND_1531 = {1{`RANDOM}};
  frameBuffer_11_107 = _RAND_1531[7:0];
  _RAND_1532 = {1{`RANDOM}};
  frameBuffer_11_108 = _RAND_1532[7:0];
  _RAND_1533 = {1{`RANDOM}};
  frameBuffer_11_109 = _RAND_1533[7:0];
  _RAND_1534 = {1{`RANDOM}};
  frameBuffer_11_110 = _RAND_1534[7:0];
  _RAND_1535 = {1{`RANDOM}};
  frameBuffer_11_111 = _RAND_1535[7:0];
  _RAND_1536 = {1{`RANDOM}};
  frameBuffer_11_112 = _RAND_1536[7:0];
  _RAND_1537 = {1{`RANDOM}};
  frameBuffer_11_113 = _RAND_1537[7:0];
  _RAND_1538 = {1{`RANDOM}};
  frameBuffer_11_114 = _RAND_1538[7:0];
  _RAND_1539 = {1{`RANDOM}};
  frameBuffer_11_115 = _RAND_1539[7:0];
  _RAND_1540 = {1{`RANDOM}};
  frameBuffer_11_116 = _RAND_1540[7:0];
  _RAND_1541 = {1{`RANDOM}};
  frameBuffer_11_117 = _RAND_1541[7:0];
  _RAND_1542 = {1{`RANDOM}};
  frameBuffer_11_118 = _RAND_1542[7:0];
  _RAND_1543 = {1{`RANDOM}};
  frameBuffer_11_119 = _RAND_1543[7:0];
  _RAND_1544 = {1{`RANDOM}};
  frameBuffer_11_120 = _RAND_1544[7:0];
  _RAND_1545 = {1{`RANDOM}};
  frameBuffer_11_121 = _RAND_1545[7:0];
  _RAND_1546 = {1{`RANDOM}};
  frameBuffer_11_122 = _RAND_1546[7:0];
  _RAND_1547 = {1{`RANDOM}};
  frameBuffer_11_123 = _RAND_1547[7:0];
  _RAND_1548 = {1{`RANDOM}};
  frameBuffer_11_124 = _RAND_1548[7:0];
  _RAND_1549 = {1{`RANDOM}};
  frameBuffer_11_125 = _RAND_1549[7:0];
  _RAND_1550 = {1{`RANDOM}};
  frameBuffer_11_126 = _RAND_1550[7:0];
  _RAND_1551 = {1{`RANDOM}};
  frameBuffer_11_127 = _RAND_1551[7:0];
  _RAND_1552 = {1{`RANDOM}};
  frameBuffer_12_0 = _RAND_1552[7:0];
  _RAND_1553 = {1{`RANDOM}};
  frameBuffer_12_1 = _RAND_1553[7:0];
  _RAND_1554 = {1{`RANDOM}};
  frameBuffer_12_2 = _RAND_1554[7:0];
  _RAND_1555 = {1{`RANDOM}};
  frameBuffer_12_3 = _RAND_1555[7:0];
  _RAND_1556 = {1{`RANDOM}};
  frameBuffer_12_4 = _RAND_1556[7:0];
  _RAND_1557 = {1{`RANDOM}};
  frameBuffer_12_5 = _RAND_1557[7:0];
  _RAND_1558 = {1{`RANDOM}};
  frameBuffer_12_6 = _RAND_1558[7:0];
  _RAND_1559 = {1{`RANDOM}};
  frameBuffer_12_7 = _RAND_1559[7:0];
  _RAND_1560 = {1{`RANDOM}};
  frameBuffer_12_8 = _RAND_1560[7:0];
  _RAND_1561 = {1{`RANDOM}};
  frameBuffer_12_9 = _RAND_1561[7:0];
  _RAND_1562 = {1{`RANDOM}};
  frameBuffer_12_10 = _RAND_1562[7:0];
  _RAND_1563 = {1{`RANDOM}};
  frameBuffer_12_11 = _RAND_1563[7:0];
  _RAND_1564 = {1{`RANDOM}};
  frameBuffer_12_12 = _RAND_1564[7:0];
  _RAND_1565 = {1{`RANDOM}};
  frameBuffer_12_13 = _RAND_1565[7:0];
  _RAND_1566 = {1{`RANDOM}};
  frameBuffer_12_14 = _RAND_1566[7:0];
  _RAND_1567 = {1{`RANDOM}};
  frameBuffer_12_15 = _RAND_1567[7:0];
  _RAND_1568 = {1{`RANDOM}};
  frameBuffer_12_16 = _RAND_1568[7:0];
  _RAND_1569 = {1{`RANDOM}};
  frameBuffer_12_17 = _RAND_1569[7:0];
  _RAND_1570 = {1{`RANDOM}};
  frameBuffer_12_18 = _RAND_1570[7:0];
  _RAND_1571 = {1{`RANDOM}};
  frameBuffer_12_19 = _RAND_1571[7:0];
  _RAND_1572 = {1{`RANDOM}};
  frameBuffer_12_20 = _RAND_1572[7:0];
  _RAND_1573 = {1{`RANDOM}};
  frameBuffer_12_21 = _RAND_1573[7:0];
  _RAND_1574 = {1{`RANDOM}};
  frameBuffer_12_22 = _RAND_1574[7:0];
  _RAND_1575 = {1{`RANDOM}};
  frameBuffer_12_23 = _RAND_1575[7:0];
  _RAND_1576 = {1{`RANDOM}};
  frameBuffer_12_24 = _RAND_1576[7:0];
  _RAND_1577 = {1{`RANDOM}};
  frameBuffer_12_25 = _RAND_1577[7:0];
  _RAND_1578 = {1{`RANDOM}};
  frameBuffer_12_26 = _RAND_1578[7:0];
  _RAND_1579 = {1{`RANDOM}};
  frameBuffer_12_27 = _RAND_1579[7:0];
  _RAND_1580 = {1{`RANDOM}};
  frameBuffer_12_28 = _RAND_1580[7:0];
  _RAND_1581 = {1{`RANDOM}};
  frameBuffer_12_29 = _RAND_1581[7:0];
  _RAND_1582 = {1{`RANDOM}};
  frameBuffer_12_30 = _RAND_1582[7:0];
  _RAND_1583 = {1{`RANDOM}};
  frameBuffer_12_31 = _RAND_1583[7:0];
  _RAND_1584 = {1{`RANDOM}};
  frameBuffer_12_32 = _RAND_1584[7:0];
  _RAND_1585 = {1{`RANDOM}};
  frameBuffer_12_33 = _RAND_1585[7:0];
  _RAND_1586 = {1{`RANDOM}};
  frameBuffer_12_34 = _RAND_1586[7:0];
  _RAND_1587 = {1{`RANDOM}};
  frameBuffer_12_35 = _RAND_1587[7:0];
  _RAND_1588 = {1{`RANDOM}};
  frameBuffer_12_36 = _RAND_1588[7:0];
  _RAND_1589 = {1{`RANDOM}};
  frameBuffer_12_37 = _RAND_1589[7:0];
  _RAND_1590 = {1{`RANDOM}};
  frameBuffer_12_38 = _RAND_1590[7:0];
  _RAND_1591 = {1{`RANDOM}};
  frameBuffer_12_39 = _RAND_1591[7:0];
  _RAND_1592 = {1{`RANDOM}};
  frameBuffer_12_40 = _RAND_1592[7:0];
  _RAND_1593 = {1{`RANDOM}};
  frameBuffer_12_41 = _RAND_1593[7:0];
  _RAND_1594 = {1{`RANDOM}};
  frameBuffer_12_42 = _RAND_1594[7:0];
  _RAND_1595 = {1{`RANDOM}};
  frameBuffer_12_43 = _RAND_1595[7:0];
  _RAND_1596 = {1{`RANDOM}};
  frameBuffer_12_44 = _RAND_1596[7:0];
  _RAND_1597 = {1{`RANDOM}};
  frameBuffer_12_45 = _RAND_1597[7:0];
  _RAND_1598 = {1{`RANDOM}};
  frameBuffer_12_46 = _RAND_1598[7:0];
  _RAND_1599 = {1{`RANDOM}};
  frameBuffer_12_47 = _RAND_1599[7:0];
  _RAND_1600 = {1{`RANDOM}};
  frameBuffer_12_48 = _RAND_1600[7:0];
  _RAND_1601 = {1{`RANDOM}};
  frameBuffer_12_49 = _RAND_1601[7:0];
  _RAND_1602 = {1{`RANDOM}};
  frameBuffer_12_50 = _RAND_1602[7:0];
  _RAND_1603 = {1{`RANDOM}};
  frameBuffer_12_51 = _RAND_1603[7:0];
  _RAND_1604 = {1{`RANDOM}};
  frameBuffer_12_52 = _RAND_1604[7:0];
  _RAND_1605 = {1{`RANDOM}};
  frameBuffer_12_53 = _RAND_1605[7:0];
  _RAND_1606 = {1{`RANDOM}};
  frameBuffer_12_54 = _RAND_1606[7:0];
  _RAND_1607 = {1{`RANDOM}};
  frameBuffer_12_55 = _RAND_1607[7:0];
  _RAND_1608 = {1{`RANDOM}};
  frameBuffer_12_56 = _RAND_1608[7:0];
  _RAND_1609 = {1{`RANDOM}};
  frameBuffer_12_57 = _RAND_1609[7:0];
  _RAND_1610 = {1{`RANDOM}};
  frameBuffer_12_58 = _RAND_1610[7:0];
  _RAND_1611 = {1{`RANDOM}};
  frameBuffer_12_59 = _RAND_1611[7:0];
  _RAND_1612 = {1{`RANDOM}};
  frameBuffer_12_60 = _RAND_1612[7:0];
  _RAND_1613 = {1{`RANDOM}};
  frameBuffer_12_61 = _RAND_1613[7:0];
  _RAND_1614 = {1{`RANDOM}};
  frameBuffer_12_62 = _RAND_1614[7:0];
  _RAND_1615 = {1{`RANDOM}};
  frameBuffer_12_63 = _RAND_1615[7:0];
  _RAND_1616 = {1{`RANDOM}};
  frameBuffer_12_64 = _RAND_1616[7:0];
  _RAND_1617 = {1{`RANDOM}};
  frameBuffer_12_65 = _RAND_1617[7:0];
  _RAND_1618 = {1{`RANDOM}};
  frameBuffer_12_66 = _RAND_1618[7:0];
  _RAND_1619 = {1{`RANDOM}};
  frameBuffer_12_67 = _RAND_1619[7:0];
  _RAND_1620 = {1{`RANDOM}};
  frameBuffer_12_68 = _RAND_1620[7:0];
  _RAND_1621 = {1{`RANDOM}};
  frameBuffer_12_69 = _RAND_1621[7:0];
  _RAND_1622 = {1{`RANDOM}};
  frameBuffer_12_70 = _RAND_1622[7:0];
  _RAND_1623 = {1{`RANDOM}};
  frameBuffer_12_71 = _RAND_1623[7:0];
  _RAND_1624 = {1{`RANDOM}};
  frameBuffer_12_72 = _RAND_1624[7:0];
  _RAND_1625 = {1{`RANDOM}};
  frameBuffer_12_73 = _RAND_1625[7:0];
  _RAND_1626 = {1{`RANDOM}};
  frameBuffer_12_74 = _RAND_1626[7:0];
  _RAND_1627 = {1{`RANDOM}};
  frameBuffer_12_75 = _RAND_1627[7:0];
  _RAND_1628 = {1{`RANDOM}};
  frameBuffer_12_76 = _RAND_1628[7:0];
  _RAND_1629 = {1{`RANDOM}};
  frameBuffer_12_77 = _RAND_1629[7:0];
  _RAND_1630 = {1{`RANDOM}};
  frameBuffer_12_78 = _RAND_1630[7:0];
  _RAND_1631 = {1{`RANDOM}};
  frameBuffer_12_79 = _RAND_1631[7:0];
  _RAND_1632 = {1{`RANDOM}};
  frameBuffer_12_80 = _RAND_1632[7:0];
  _RAND_1633 = {1{`RANDOM}};
  frameBuffer_12_81 = _RAND_1633[7:0];
  _RAND_1634 = {1{`RANDOM}};
  frameBuffer_12_82 = _RAND_1634[7:0];
  _RAND_1635 = {1{`RANDOM}};
  frameBuffer_12_83 = _RAND_1635[7:0];
  _RAND_1636 = {1{`RANDOM}};
  frameBuffer_12_84 = _RAND_1636[7:0];
  _RAND_1637 = {1{`RANDOM}};
  frameBuffer_12_85 = _RAND_1637[7:0];
  _RAND_1638 = {1{`RANDOM}};
  frameBuffer_12_86 = _RAND_1638[7:0];
  _RAND_1639 = {1{`RANDOM}};
  frameBuffer_12_87 = _RAND_1639[7:0];
  _RAND_1640 = {1{`RANDOM}};
  frameBuffer_12_88 = _RAND_1640[7:0];
  _RAND_1641 = {1{`RANDOM}};
  frameBuffer_12_89 = _RAND_1641[7:0];
  _RAND_1642 = {1{`RANDOM}};
  frameBuffer_12_90 = _RAND_1642[7:0];
  _RAND_1643 = {1{`RANDOM}};
  frameBuffer_12_91 = _RAND_1643[7:0];
  _RAND_1644 = {1{`RANDOM}};
  frameBuffer_12_92 = _RAND_1644[7:0];
  _RAND_1645 = {1{`RANDOM}};
  frameBuffer_12_93 = _RAND_1645[7:0];
  _RAND_1646 = {1{`RANDOM}};
  frameBuffer_12_94 = _RAND_1646[7:0];
  _RAND_1647 = {1{`RANDOM}};
  frameBuffer_12_95 = _RAND_1647[7:0];
  _RAND_1648 = {1{`RANDOM}};
  frameBuffer_12_96 = _RAND_1648[7:0];
  _RAND_1649 = {1{`RANDOM}};
  frameBuffer_12_97 = _RAND_1649[7:0];
  _RAND_1650 = {1{`RANDOM}};
  frameBuffer_12_98 = _RAND_1650[7:0];
  _RAND_1651 = {1{`RANDOM}};
  frameBuffer_12_99 = _RAND_1651[7:0];
  _RAND_1652 = {1{`RANDOM}};
  frameBuffer_12_100 = _RAND_1652[7:0];
  _RAND_1653 = {1{`RANDOM}};
  frameBuffer_12_101 = _RAND_1653[7:0];
  _RAND_1654 = {1{`RANDOM}};
  frameBuffer_12_102 = _RAND_1654[7:0];
  _RAND_1655 = {1{`RANDOM}};
  frameBuffer_12_103 = _RAND_1655[7:0];
  _RAND_1656 = {1{`RANDOM}};
  frameBuffer_12_104 = _RAND_1656[7:0];
  _RAND_1657 = {1{`RANDOM}};
  frameBuffer_12_105 = _RAND_1657[7:0];
  _RAND_1658 = {1{`RANDOM}};
  frameBuffer_12_106 = _RAND_1658[7:0];
  _RAND_1659 = {1{`RANDOM}};
  frameBuffer_12_107 = _RAND_1659[7:0];
  _RAND_1660 = {1{`RANDOM}};
  frameBuffer_12_108 = _RAND_1660[7:0];
  _RAND_1661 = {1{`RANDOM}};
  frameBuffer_12_109 = _RAND_1661[7:0];
  _RAND_1662 = {1{`RANDOM}};
  frameBuffer_12_110 = _RAND_1662[7:0];
  _RAND_1663 = {1{`RANDOM}};
  frameBuffer_12_111 = _RAND_1663[7:0];
  _RAND_1664 = {1{`RANDOM}};
  frameBuffer_12_112 = _RAND_1664[7:0];
  _RAND_1665 = {1{`RANDOM}};
  frameBuffer_12_113 = _RAND_1665[7:0];
  _RAND_1666 = {1{`RANDOM}};
  frameBuffer_12_114 = _RAND_1666[7:0];
  _RAND_1667 = {1{`RANDOM}};
  frameBuffer_12_115 = _RAND_1667[7:0];
  _RAND_1668 = {1{`RANDOM}};
  frameBuffer_12_116 = _RAND_1668[7:0];
  _RAND_1669 = {1{`RANDOM}};
  frameBuffer_12_117 = _RAND_1669[7:0];
  _RAND_1670 = {1{`RANDOM}};
  frameBuffer_12_118 = _RAND_1670[7:0];
  _RAND_1671 = {1{`RANDOM}};
  frameBuffer_12_119 = _RAND_1671[7:0];
  _RAND_1672 = {1{`RANDOM}};
  frameBuffer_12_120 = _RAND_1672[7:0];
  _RAND_1673 = {1{`RANDOM}};
  frameBuffer_12_121 = _RAND_1673[7:0];
  _RAND_1674 = {1{`RANDOM}};
  frameBuffer_12_122 = _RAND_1674[7:0];
  _RAND_1675 = {1{`RANDOM}};
  frameBuffer_12_123 = _RAND_1675[7:0];
  _RAND_1676 = {1{`RANDOM}};
  frameBuffer_12_124 = _RAND_1676[7:0];
  _RAND_1677 = {1{`RANDOM}};
  frameBuffer_12_125 = _RAND_1677[7:0];
  _RAND_1678 = {1{`RANDOM}};
  frameBuffer_12_126 = _RAND_1678[7:0];
  _RAND_1679 = {1{`RANDOM}};
  frameBuffer_12_127 = _RAND_1679[7:0];
  _RAND_1680 = {1{`RANDOM}};
  frameBuffer_13_0 = _RAND_1680[7:0];
  _RAND_1681 = {1{`RANDOM}};
  frameBuffer_13_1 = _RAND_1681[7:0];
  _RAND_1682 = {1{`RANDOM}};
  frameBuffer_13_2 = _RAND_1682[7:0];
  _RAND_1683 = {1{`RANDOM}};
  frameBuffer_13_3 = _RAND_1683[7:0];
  _RAND_1684 = {1{`RANDOM}};
  frameBuffer_13_4 = _RAND_1684[7:0];
  _RAND_1685 = {1{`RANDOM}};
  frameBuffer_13_5 = _RAND_1685[7:0];
  _RAND_1686 = {1{`RANDOM}};
  frameBuffer_13_6 = _RAND_1686[7:0];
  _RAND_1687 = {1{`RANDOM}};
  frameBuffer_13_7 = _RAND_1687[7:0];
  _RAND_1688 = {1{`RANDOM}};
  frameBuffer_13_8 = _RAND_1688[7:0];
  _RAND_1689 = {1{`RANDOM}};
  frameBuffer_13_9 = _RAND_1689[7:0];
  _RAND_1690 = {1{`RANDOM}};
  frameBuffer_13_10 = _RAND_1690[7:0];
  _RAND_1691 = {1{`RANDOM}};
  frameBuffer_13_11 = _RAND_1691[7:0];
  _RAND_1692 = {1{`RANDOM}};
  frameBuffer_13_12 = _RAND_1692[7:0];
  _RAND_1693 = {1{`RANDOM}};
  frameBuffer_13_13 = _RAND_1693[7:0];
  _RAND_1694 = {1{`RANDOM}};
  frameBuffer_13_14 = _RAND_1694[7:0];
  _RAND_1695 = {1{`RANDOM}};
  frameBuffer_13_15 = _RAND_1695[7:0];
  _RAND_1696 = {1{`RANDOM}};
  frameBuffer_13_16 = _RAND_1696[7:0];
  _RAND_1697 = {1{`RANDOM}};
  frameBuffer_13_17 = _RAND_1697[7:0];
  _RAND_1698 = {1{`RANDOM}};
  frameBuffer_13_18 = _RAND_1698[7:0];
  _RAND_1699 = {1{`RANDOM}};
  frameBuffer_13_19 = _RAND_1699[7:0];
  _RAND_1700 = {1{`RANDOM}};
  frameBuffer_13_20 = _RAND_1700[7:0];
  _RAND_1701 = {1{`RANDOM}};
  frameBuffer_13_21 = _RAND_1701[7:0];
  _RAND_1702 = {1{`RANDOM}};
  frameBuffer_13_22 = _RAND_1702[7:0];
  _RAND_1703 = {1{`RANDOM}};
  frameBuffer_13_23 = _RAND_1703[7:0];
  _RAND_1704 = {1{`RANDOM}};
  frameBuffer_13_24 = _RAND_1704[7:0];
  _RAND_1705 = {1{`RANDOM}};
  frameBuffer_13_25 = _RAND_1705[7:0];
  _RAND_1706 = {1{`RANDOM}};
  frameBuffer_13_26 = _RAND_1706[7:0];
  _RAND_1707 = {1{`RANDOM}};
  frameBuffer_13_27 = _RAND_1707[7:0];
  _RAND_1708 = {1{`RANDOM}};
  frameBuffer_13_28 = _RAND_1708[7:0];
  _RAND_1709 = {1{`RANDOM}};
  frameBuffer_13_29 = _RAND_1709[7:0];
  _RAND_1710 = {1{`RANDOM}};
  frameBuffer_13_30 = _RAND_1710[7:0];
  _RAND_1711 = {1{`RANDOM}};
  frameBuffer_13_31 = _RAND_1711[7:0];
  _RAND_1712 = {1{`RANDOM}};
  frameBuffer_13_32 = _RAND_1712[7:0];
  _RAND_1713 = {1{`RANDOM}};
  frameBuffer_13_33 = _RAND_1713[7:0];
  _RAND_1714 = {1{`RANDOM}};
  frameBuffer_13_34 = _RAND_1714[7:0];
  _RAND_1715 = {1{`RANDOM}};
  frameBuffer_13_35 = _RAND_1715[7:0];
  _RAND_1716 = {1{`RANDOM}};
  frameBuffer_13_36 = _RAND_1716[7:0];
  _RAND_1717 = {1{`RANDOM}};
  frameBuffer_13_37 = _RAND_1717[7:0];
  _RAND_1718 = {1{`RANDOM}};
  frameBuffer_13_38 = _RAND_1718[7:0];
  _RAND_1719 = {1{`RANDOM}};
  frameBuffer_13_39 = _RAND_1719[7:0];
  _RAND_1720 = {1{`RANDOM}};
  frameBuffer_13_40 = _RAND_1720[7:0];
  _RAND_1721 = {1{`RANDOM}};
  frameBuffer_13_41 = _RAND_1721[7:0];
  _RAND_1722 = {1{`RANDOM}};
  frameBuffer_13_42 = _RAND_1722[7:0];
  _RAND_1723 = {1{`RANDOM}};
  frameBuffer_13_43 = _RAND_1723[7:0];
  _RAND_1724 = {1{`RANDOM}};
  frameBuffer_13_44 = _RAND_1724[7:0];
  _RAND_1725 = {1{`RANDOM}};
  frameBuffer_13_45 = _RAND_1725[7:0];
  _RAND_1726 = {1{`RANDOM}};
  frameBuffer_13_46 = _RAND_1726[7:0];
  _RAND_1727 = {1{`RANDOM}};
  frameBuffer_13_47 = _RAND_1727[7:0];
  _RAND_1728 = {1{`RANDOM}};
  frameBuffer_13_48 = _RAND_1728[7:0];
  _RAND_1729 = {1{`RANDOM}};
  frameBuffer_13_49 = _RAND_1729[7:0];
  _RAND_1730 = {1{`RANDOM}};
  frameBuffer_13_50 = _RAND_1730[7:0];
  _RAND_1731 = {1{`RANDOM}};
  frameBuffer_13_51 = _RAND_1731[7:0];
  _RAND_1732 = {1{`RANDOM}};
  frameBuffer_13_52 = _RAND_1732[7:0];
  _RAND_1733 = {1{`RANDOM}};
  frameBuffer_13_53 = _RAND_1733[7:0];
  _RAND_1734 = {1{`RANDOM}};
  frameBuffer_13_54 = _RAND_1734[7:0];
  _RAND_1735 = {1{`RANDOM}};
  frameBuffer_13_55 = _RAND_1735[7:0];
  _RAND_1736 = {1{`RANDOM}};
  frameBuffer_13_56 = _RAND_1736[7:0];
  _RAND_1737 = {1{`RANDOM}};
  frameBuffer_13_57 = _RAND_1737[7:0];
  _RAND_1738 = {1{`RANDOM}};
  frameBuffer_13_58 = _RAND_1738[7:0];
  _RAND_1739 = {1{`RANDOM}};
  frameBuffer_13_59 = _RAND_1739[7:0];
  _RAND_1740 = {1{`RANDOM}};
  frameBuffer_13_60 = _RAND_1740[7:0];
  _RAND_1741 = {1{`RANDOM}};
  frameBuffer_13_61 = _RAND_1741[7:0];
  _RAND_1742 = {1{`RANDOM}};
  frameBuffer_13_62 = _RAND_1742[7:0];
  _RAND_1743 = {1{`RANDOM}};
  frameBuffer_13_63 = _RAND_1743[7:0];
  _RAND_1744 = {1{`RANDOM}};
  frameBuffer_13_64 = _RAND_1744[7:0];
  _RAND_1745 = {1{`RANDOM}};
  frameBuffer_13_65 = _RAND_1745[7:0];
  _RAND_1746 = {1{`RANDOM}};
  frameBuffer_13_66 = _RAND_1746[7:0];
  _RAND_1747 = {1{`RANDOM}};
  frameBuffer_13_67 = _RAND_1747[7:0];
  _RAND_1748 = {1{`RANDOM}};
  frameBuffer_13_68 = _RAND_1748[7:0];
  _RAND_1749 = {1{`RANDOM}};
  frameBuffer_13_69 = _RAND_1749[7:0];
  _RAND_1750 = {1{`RANDOM}};
  frameBuffer_13_70 = _RAND_1750[7:0];
  _RAND_1751 = {1{`RANDOM}};
  frameBuffer_13_71 = _RAND_1751[7:0];
  _RAND_1752 = {1{`RANDOM}};
  frameBuffer_13_72 = _RAND_1752[7:0];
  _RAND_1753 = {1{`RANDOM}};
  frameBuffer_13_73 = _RAND_1753[7:0];
  _RAND_1754 = {1{`RANDOM}};
  frameBuffer_13_74 = _RAND_1754[7:0];
  _RAND_1755 = {1{`RANDOM}};
  frameBuffer_13_75 = _RAND_1755[7:0];
  _RAND_1756 = {1{`RANDOM}};
  frameBuffer_13_76 = _RAND_1756[7:0];
  _RAND_1757 = {1{`RANDOM}};
  frameBuffer_13_77 = _RAND_1757[7:0];
  _RAND_1758 = {1{`RANDOM}};
  frameBuffer_13_78 = _RAND_1758[7:0];
  _RAND_1759 = {1{`RANDOM}};
  frameBuffer_13_79 = _RAND_1759[7:0];
  _RAND_1760 = {1{`RANDOM}};
  frameBuffer_13_80 = _RAND_1760[7:0];
  _RAND_1761 = {1{`RANDOM}};
  frameBuffer_13_81 = _RAND_1761[7:0];
  _RAND_1762 = {1{`RANDOM}};
  frameBuffer_13_82 = _RAND_1762[7:0];
  _RAND_1763 = {1{`RANDOM}};
  frameBuffer_13_83 = _RAND_1763[7:0];
  _RAND_1764 = {1{`RANDOM}};
  frameBuffer_13_84 = _RAND_1764[7:0];
  _RAND_1765 = {1{`RANDOM}};
  frameBuffer_13_85 = _RAND_1765[7:0];
  _RAND_1766 = {1{`RANDOM}};
  frameBuffer_13_86 = _RAND_1766[7:0];
  _RAND_1767 = {1{`RANDOM}};
  frameBuffer_13_87 = _RAND_1767[7:0];
  _RAND_1768 = {1{`RANDOM}};
  frameBuffer_13_88 = _RAND_1768[7:0];
  _RAND_1769 = {1{`RANDOM}};
  frameBuffer_13_89 = _RAND_1769[7:0];
  _RAND_1770 = {1{`RANDOM}};
  frameBuffer_13_90 = _RAND_1770[7:0];
  _RAND_1771 = {1{`RANDOM}};
  frameBuffer_13_91 = _RAND_1771[7:0];
  _RAND_1772 = {1{`RANDOM}};
  frameBuffer_13_92 = _RAND_1772[7:0];
  _RAND_1773 = {1{`RANDOM}};
  frameBuffer_13_93 = _RAND_1773[7:0];
  _RAND_1774 = {1{`RANDOM}};
  frameBuffer_13_94 = _RAND_1774[7:0];
  _RAND_1775 = {1{`RANDOM}};
  frameBuffer_13_95 = _RAND_1775[7:0];
  _RAND_1776 = {1{`RANDOM}};
  frameBuffer_13_96 = _RAND_1776[7:0];
  _RAND_1777 = {1{`RANDOM}};
  frameBuffer_13_97 = _RAND_1777[7:0];
  _RAND_1778 = {1{`RANDOM}};
  frameBuffer_13_98 = _RAND_1778[7:0];
  _RAND_1779 = {1{`RANDOM}};
  frameBuffer_13_99 = _RAND_1779[7:0];
  _RAND_1780 = {1{`RANDOM}};
  frameBuffer_13_100 = _RAND_1780[7:0];
  _RAND_1781 = {1{`RANDOM}};
  frameBuffer_13_101 = _RAND_1781[7:0];
  _RAND_1782 = {1{`RANDOM}};
  frameBuffer_13_102 = _RAND_1782[7:0];
  _RAND_1783 = {1{`RANDOM}};
  frameBuffer_13_103 = _RAND_1783[7:0];
  _RAND_1784 = {1{`RANDOM}};
  frameBuffer_13_104 = _RAND_1784[7:0];
  _RAND_1785 = {1{`RANDOM}};
  frameBuffer_13_105 = _RAND_1785[7:0];
  _RAND_1786 = {1{`RANDOM}};
  frameBuffer_13_106 = _RAND_1786[7:0];
  _RAND_1787 = {1{`RANDOM}};
  frameBuffer_13_107 = _RAND_1787[7:0];
  _RAND_1788 = {1{`RANDOM}};
  frameBuffer_13_108 = _RAND_1788[7:0];
  _RAND_1789 = {1{`RANDOM}};
  frameBuffer_13_109 = _RAND_1789[7:0];
  _RAND_1790 = {1{`RANDOM}};
  frameBuffer_13_110 = _RAND_1790[7:0];
  _RAND_1791 = {1{`RANDOM}};
  frameBuffer_13_111 = _RAND_1791[7:0];
  _RAND_1792 = {1{`RANDOM}};
  frameBuffer_13_112 = _RAND_1792[7:0];
  _RAND_1793 = {1{`RANDOM}};
  frameBuffer_13_113 = _RAND_1793[7:0];
  _RAND_1794 = {1{`RANDOM}};
  frameBuffer_13_114 = _RAND_1794[7:0];
  _RAND_1795 = {1{`RANDOM}};
  frameBuffer_13_115 = _RAND_1795[7:0];
  _RAND_1796 = {1{`RANDOM}};
  frameBuffer_13_116 = _RAND_1796[7:0];
  _RAND_1797 = {1{`RANDOM}};
  frameBuffer_13_117 = _RAND_1797[7:0];
  _RAND_1798 = {1{`RANDOM}};
  frameBuffer_13_118 = _RAND_1798[7:0];
  _RAND_1799 = {1{`RANDOM}};
  frameBuffer_13_119 = _RAND_1799[7:0];
  _RAND_1800 = {1{`RANDOM}};
  frameBuffer_13_120 = _RAND_1800[7:0];
  _RAND_1801 = {1{`RANDOM}};
  frameBuffer_13_121 = _RAND_1801[7:0];
  _RAND_1802 = {1{`RANDOM}};
  frameBuffer_13_122 = _RAND_1802[7:0];
  _RAND_1803 = {1{`RANDOM}};
  frameBuffer_13_123 = _RAND_1803[7:0];
  _RAND_1804 = {1{`RANDOM}};
  frameBuffer_13_124 = _RAND_1804[7:0];
  _RAND_1805 = {1{`RANDOM}};
  frameBuffer_13_125 = _RAND_1805[7:0];
  _RAND_1806 = {1{`RANDOM}};
  frameBuffer_13_126 = _RAND_1806[7:0];
  _RAND_1807 = {1{`RANDOM}};
  frameBuffer_13_127 = _RAND_1807[7:0];
  _RAND_1808 = {1{`RANDOM}};
  frameBuffer_14_0 = _RAND_1808[7:0];
  _RAND_1809 = {1{`RANDOM}};
  frameBuffer_14_1 = _RAND_1809[7:0];
  _RAND_1810 = {1{`RANDOM}};
  frameBuffer_14_2 = _RAND_1810[7:0];
  _RAND_1811 = {1{`RANDOM}};
  frameBuffer_14_3 = _RAND_1811[7:0];
  _RAND_1812 = {1{`RANDOM}};
  frameBuffer_14_4 = _RAND_1812[7:0];
  _RAND_1813 = {1{`RANDOM}};
  frameBuffer_14_5 = _RAND_1813[7:0];
  _RAND_1814 = {1{`RANDOM}};
  frameBuffer_14_6 = _RAND_1814[7:0];
  _RAND_1815 = {1{`RANDOM}};
  frameBuffer_14_7 = _RAND_1815[7:0];
  _RAND_1816 = {1{`RANDOM}};
  frameBuffer_14_8 = _RAND_1816[7:0];
  _RAND_1817 = {1{`RANDOM}};
  frameBuffer_14_9 = _RAND_1817[7:0];
  _RAND_1818 = {1{`RANDOM}};
  frameBuffer_14_10 = _RAND_1818[7:0];
  _RAND_1819 = {1{`RANDOM}};
  frameBuffer_14_11 = _RAND_1819[7:0];
  _RAND_1820 = {1{`RANDOM}};
  frameBuffer_14_12 = _RAND_1820[7:0];
  _RAND_1821 = {1{`RANDOM}};
  frameBuffer_14_13 = _RAND_1821[7:0];
  _RAND_1822 = {1{`RANDOM}};
  frameBuffer_14_14 = _RAND_1822[7:0];
  _RAND_1823 = {1{`RANDOM}};
  frameBuffer_14_15 = _RAND_1823[7:0];
  _RAND_1824 = {1{`RANDOM}};
  frameBuffer_14_16 = _RAND_1824[7:0];
  _RAND_1825 = {1{`RANDOM}};
  frameBuffer_14_17 = _RAND_1825[7:0];
  _RAND_1826 = {1{`RANDOM}};
  frameBuffer_14_18 = _RAND_1826[7:0];
  _RAND_1827 = {1{`RANDOM}};
  frameBuffer_14_19 = _RAND_1827[7:0];
  _RAND_1828 = {1{`RANDOM}};
  frameBuffer_14_20 = _RAND_1828[7:0];
  _RAND_1829 = {1{`RANDOM}};
  frameBuffer_14_21 = _RAND_1829[7:0];
  _RAND_1830 = {1{`RANDOM}};
  frameBuffer_14_22 = _RAND_1830[7:0];
  _RAND_1831 = {1{`RANDOM}};
  frameBuffer_14_23 = _RAND_1831[7:0];
  _RAND_1832 = {1{`RANDOM}};
  frameBuffer_14_24 = _RAND_1832[7:0];
  _RAND_1833 = {1{`RANDOM}};
  frameBuffer_14_25 = _RAND_1833[7:0];
  _RAND_1834 = {1{`RANDOM}};
  frameBuffer_14_26 = _RAND_1834[7:0];
  _RAND_1835 = {1{`RANDOM}};
  frameBuffer_14_27 = _RAND_1835[7:0];
  _RAND_1836 = {1{`RANDOM}};
  frameBuffer_14_28 = _RAND_1836[7:0];
  _RAND_1837 = {1{`RANDOM}};
  frameBuffer_14_29 = _RAND_1837[7:0];
  _RAND_1838 = {1{`RANDOM}};
  frameBuffer_14_30 = _RAND_1838[7:0];
  _RAND_1839 = {1{`RANDOM}};
  frameBuffer_14_31 = _RAND_1839[7:0];
  _RAND_1840 = {1{`RANDOM}};
  frameBuffer_14_32 = _RAND_1840[7:0];
  _RAND_1841 = {1{`RANDOM}};
  frameBuffer_14_33 = _RAND_1841[7:0];
  _RAND_1842 = {1{`RANDOM}};
  frameBuffer_14_34 = _RAND_1842[7:0];
  _RAND_1843 = {1{`RANDOM}};
  frameBuffer_14_35 = _RAND_1843[7:0];
  _RAND_1844 = {1{`RANDOM}};
  frameBuffer_14_36 = _RAND_1844[7:0];
  _RAND_1845 = {1{`RANDOM}};
  frameBuffer_14_37 = _RAND_1845[7:0];
  _RAND_1846 = {1{`RANDOM}};
  frameBuffer_14_38 = _RAND_1846[7:0];
  _RAND_1847 = {1{`RANDOM}};
  frameBuffer_14_39 = _RAND_1847[7:0];
  _RAND_1848 = {1{`RANDOM}};
  frameBuffer_14_40 = _RAND_1848[7:0];
  _RAND_1849 = {1{`RANDOM}};
  frameBuffer_14_41 = _RAND_1849[7:0];
  _RAND_1850 = {1{`RANDOM}};
  frameBuffer_14_42 = _RAND_1850[7:0];
  _RAND_1851 = {1{`RANDOM}};
  frameBuffer_14_43 = _RAND_1851[7:0];
  _RAND_1852 = {1{`RANDOM}};
  frameBuffer_14_44 = _RAND_1852[7:0];
  _RAND_1853 = {1{`RANDOM}};
  frameBuffer_14_45 = _RAND_1853[7:0];
  _RAND_1854 = {1{`RANDOM}};
  frameBuffer_14_46 = _RAND_1854[7:0];
  _RAND_1855 = {1{`RANDOM}};
  frameBuffer_14_47 = _RAND_1855[7:0];
  _RAND_1856 = {1{`RANDOM}};
  frameBuffer_14_48 = _RAND_1856[7:0];
  _RAND_1857 = {1{`RANDOM}};
  frameBuffer_14_49 = _RAND_1857[7:0];
  _RAND_1858 = {1{`RANDOM}};
  frameBuffer_14_50 = _RAND_1858[7:0];
  _RAND_1859 = {1{`RANDOM}};
  frameBuffer_14_51 = _RAND_1859[7:0];
  _RAND_1860 = {1{`RANDOM}};
  frameBuffer_14_52 = _RAND_1860[7:0];
  _RAND_1861 = {1{`RANDOM}};
  frameBuffer_14_53 = _RAND_1861[7:0];
  _RAND_1862 = {1{`RANDOM}};
  frameBuffer_14_54 = _RAND_1862[7:0];
  _RAND_1863 = {1{`RANDOM}};
  frameBuffer_14_55 = _RAND_1863[7:0];
  _RAND_1864 = {1{`RANDOM}};
  frameBuffer_14_56 = _RAND_1864[7:0];
  _RAND_1865 = {1{`RANDOM}};
  frameBuffer_14_57 = _RAND_1865[7:0];
  _RAND_1866 = {1{`RANDOM}};
  frameBuffer_14_58 = _RAND_1866[7:0];
  _RAND_1867 = {1{`RANDOM}};
  frameBuffer_14_59 = _RAND_1867[7:0];
  _RAND_1868 = {1{`RANDOM}};
  frameBuffer_14_60 = _RAND_1868[7:0];
  _RAND_1869 = {1{`RANDOM}};
  frameBuffer_14_61 = _RAND_1869[7:0];
  _RAND_1870 = {1{`RANDOM}};
  frameBuffer_14_62 = _RAND_1870[7:0];
  _RAND_1871 = {1{`RANDOM}};
  frameBuffer_14_63 = _RAND_1871[7:0];
  _RAND_1872 = {1{`RANDOM}};
  frameBuffer_14_64 = _RAND_1872[7:0];
  _RAND_1873 = {1{`RANDOM}};
  frameBuffer_14_65 = _RAND_1873[7:0];
  _RAND_1874 = {1{`RANDOM}};
  frameBuffer_14_66 = _RAND_1874[7:0];
  _RAND_1875 = {1{`RANDOM}};
  frameBuffer_14_67 = _RAND_1875[7:0];
  _RAND_1876 = {1{`RANDOM}};
  frameBuffer_14_68 = _RAND_1876[7:0];
  _RAND_1877 = {1{`RANDOM}};
  frameBuffer_14_69 = _RAND_1877[7:0];
  _RAND_1878 = {1{`RANDOM}};
  frameBuffer_14_70 = _RAND_1878[7:0];
  _RAND_1879 = {1{`RANDOM}};
  frameBuffer_14_71 = _RAND_1879[7:0];
  _RAND_1880 = {1{`RANDOM}};
  frameBuffer_14_72 = _RAND_1880[7:0];
  _RAND_1881 = {1{`RANDOM}};
  frameBuffer_14_73 = _RAND_1881[7:0];
  _RAND_1882 = {1{`RANDOM}};
  frameBuffer_14_74 = _RAND_1882[7:0];
  _RAND_1883 = {1{`RANDOM}};
  frameBuffer_14_75 = _RAND_1883[7:0];
  _RAND_1884 = {1{`RANDOM}};
  frameBuffer_14_76 = _RAND_1884[7:0];
  _RAND_1885 = {1{`RANDOM}};
  frameBuffer_14_77 = _RAND_1885[7:0];
  _RAND_1886 = {1{`RANDOM}};
  frameBuffer_14_78 = _RAND_1886[7:0];
  _RAND_1887 = {1{`RANDOM}};
  frameBuffer_14_79 = _RAND_1887[7:0];
  _RAND_1888 = {1{`RANDOM}};
  frameBuffer_14_80 = _RAND_1888[7:0];
  _RAND_1889 = {1{`RANDOM}};
  frameBuffer_14_81 = _RAND_1889[7:0];
  _RAND_1890 = {1{`RANDOM}};
  frameBuffer_14_82 = _RAND_1890[7:0];
  _RAND_1891 = {1{`RANDOM}};
  frameBuffer_14_83 = _RAND_1891[7:0];
  _RAND_1892 = {1{`RANDOM}};
  frameBuffer_14_84 = _RAND_1892[7:0];
  _RAND_1893 = {1{`RANDOM}};
  frameBuffer_14_85 = _RAND_1893[7:0];
  _RAND_1894 = {1{`RANDOM}};
  frameBuffer_14_86 = _RAND_1894[7:0];
  _RAND_1895 = {1{`RANDOM}};
  frameBuffer_14_87 = _RAND_1895[7:0];
  _RAND_1896 = {1{`RANDOM}};
  frameBuffer_14_88 = _RAND_1896[7:0];
  _RAND_1897 = {1{`RANDOM}};
  frameBuffer_14_89 = _RAND_1897[7:0];
  _RAND_1898 = {1{`RANDOM}};
  frameBuffer_14_90 = _RAND_1898[7:0];
  _RAND_1899 = {1{`RANDOM}};
  frameBuffer_14_91 = _RAND_1899[7:0];
  _RAND_1900 = {1{`RANDOM}};
  frameBuffer_14_92 = _RAND_1900[7:0];
  _RAND_1901 = {1{`RANDOM}};
  frameBuffer_14_93 = _RAND_1901[7:0];
  _RAND_1902 = {1{`RANDOM}};
  frameBuffer_14_94 = _RAND_1902[7:0];
  _RAND_1903 = {1{`RANDOM}};
  frameBuffer_14_95 = _RAND_1903[7:0];
  _RAND_1904 = {1{`RANDOM}};
  frameBuffer_14_96 = _RAND_1904[7:0];
  _RAND_1905 = {1{`RANDOM}};
  frameBuffer_14_97 = _RAND_1905[7:0];
  _RAND_1906 = {1{`RANDOM}};
  frameBuffer_14_98 = _RAND_1906[7:0];
  _RAND_1907 = {1{`RANDOM}};
  frameBuffer_14_99 = _RAND_1907[7:0];
  _RAND_1908 = {1{`RANDOM}};
  frameBuffer_14_100 = _RAND_1908[7:0];
  _RAND_1909 = {1{`RANDOM}};
  frameBuffer_14_101 = _RAND_1909[7:0];
  _RAND_1910 = {1{`RANDOM}};
  frameBuffer_14_102 = _RAND_1910[7:0];
  _RAND_1911 = {1{`RANDOM}};
  frameBuffer_14_103 = _RAND_1911[7:0];
  _RAND_1912 = {1{`RANDOM}};
  frameBuffer_14_104 = _RAND_1912[7:0];
  _RAND_1913 = {1{`RANDOM}};
  frameBuffer_14_105 = _RAND_1913[7:0];
  _RAND_1914 = {1{`RANDOM}};
  frameBuffer_14_106 = _RAND_1914[7:0];
  _RAND_1915 = {1{`RANDOM}};
  frameBuffer_14_107 = _RAND_1915[7:0];
  _RAND_1916 = {1{`RANDOM}};
  frameBuffer_14_108 = _RAND_1916[7:0];
  _RAND_1917 = {1{`RANDOM}};
  frameBuffer_14_109 = _RAND_1917[7:0];
  _RAND_1918 = {1{`RANDOM}};
  frameBuffer_14_110 = _RAND_1918[7:0];
  _RAND_1919 = {1{`RANDOM}};
  frameBuffer_14_111 = _RAND_1919[7:0];
  _RAND_1920 = {1{`RANDOM}};
  frameBuffer_14_112 = _RAND_1920[7:0];
  _RAND_1921 = {1{`RANDOM}};
  frameBuffer_14_113 = _RAND_1921[7:0];
  _RAND_1922 = {1{`RANDOM}};
  frameBuffer_14_114 = _RAND_1922[7:0];
  _RAND_1923 = {1{`RANDOM}};
  frameBuffer_14_115 = _RAND_1923[7:0];
  _RAND_1924 = {1{`RANDOM}};
  frameBuffer_14_116 = _RAND_1924[7:0];
  _RAND_1925 = {1{`RANDOM}};
  frameBuffer_14_117 = _RAND_1925[7:0];
  _RAND_1926 = {1{`RANDOM}};
  frameBuffer_14_118 = _RAND_1926[7:0];
  _RAND_1927 = {1{`RANDOM}};
  frameBuffer_14_119 = _RAND_1927[7:0];
  _RAND_1928 = {1{`RANDOM}};
  frameBuffer_14_120 = _RAND_1928[7:0];
  _RAND_1929 = {1{`RANDOM}};
  frameBuffer_14_121 = _RAND_1929[7:0];
  _RAND_1930 = {1{`RANDOM}};
  frameBuffer_14_122 = _RAND_1930[7:0];
  _RAND_1931 = {1{`RANDOM}};
  frameBuffer_14_123 = _RAND_1931[7:0];
  _RAND_1932 = {1{`RANDOM}};
  frameBuffer_14_124 = _RAND_1932[7:0];
  _RAND_1933 = {1{`RANDOM}};
  frameBuffer_14_125 = _RAND_1933[7:0];
  _RAND_1934 = {1{`RANDOM}};
  frameBuffer_14_126 = _RAND_1934[7:0];
  _RAND_1935 = {1{`RANDOM}};
  frameBuffer_14_127 = _RAND_1935[7:0];
  _RAND_1936 = {1{`RANDOM}};
  frameBuffer_15_0 = _RAND_1936[7:0];
  _RAND_1937 = {1{`RANDOM}};
  frameBuffer_15_1 = _RAND_1937[7:0];
  _RAND_1938 = {1{`RANDOM}};
  frameBuffer_15_2 = _RAND_1938[7:0];
  _RAND_1939 = {1{`RANDOM}};
  frameBuffer_15_3 = _RAND_1939[7:0];
  _RAND_1940 = {1{`RANDOM}};
  frameBuffer_15_4 = _RAND_1940[7:0];
  _RAND_1941 = {1{`RANDOM}};
  frameBuffer_15_5 = _RAND_1941[7:0];
  _RAND_1942 = {1{`RANDOM}};
  frameBuffer_15_6 = _RAND_1942[7:0];
  _RAND_1943 = {1{`RANDOM}};
  frameBuffer_15_7 = _RAND_1943[7:0];
  _RAND_1944 = {1{`RANDOM}};
  frameBuffer_15_8 = _RAND_1944[7:0];
  _RAND_1945 = {1{`RANDOM}};
  frameBuffer_15_9 = _RAND_1945[7:0];
  _RAND_1946 = {1{`RANDOM}};
  frameBuffer_15_10 = _RAND_1946[7:0];
  _RAND_1947 = {1{`RANDOM}};
  frameBuffer_15_11 = _RAND_1947[7:0];
  _RAND_1948 = {1{`RANDOM}};
  frameBuffer_15_12 = _RAND_1948[7:0];
  _RAND_1949 = {1{`RANDOM}};
  frameBuffer_15_13 = _RAND_1949[7:0];
  _RAND_1950 = {1{`RANDOM}};
  frameBuffer_15_14 = _RAND_1950[7:0];
  _RAND_1951 = {1{`RANDOM}};
  frameBuffer_15_15 = _RAND_1951[7:0];
  _RAND_1952 = {1{`RANDOM}};
  frameBuffer_15_16 = _RAND_1952[7:0];
  _RAND_1953 = {1{`RANDOM}};
  frameBuffer_15_17 = _RAND_1953[7:0];
  _RAND_1954 = {1{`RANDOM}};
  frameBuffer_15_18 = _RAND_1954[7:0];
  _RAND_1955 = {1{`RANDOM}};
  frameBuffer_15_19 = _RAND_1955[7:0];
  _RAND_1956 = {1{`RANDOM}};
  frameBuffer_15_20 = _RAND_1956[7:0];
  _RAND_1957 = {1{`RANDOM}};
  frameBuffer_15_21 = _RAND_1957[7:0];
  _RAND_1958 = {1{`RANDOM}};
  frameBuffer_15_22 = _RAND_1958[7:0];
  _RAND_1959 = {1{`RANDOM}};
  frameBuffer_15_23 = _RAND_1959[7:0];
  _RAND_1960 = {1{`RANDOM}};
  frameBuffer_15_24 = _RAND_1960[7:0];
  _RAND_1961 = {1{`RANDOM}};
  frameBuffer_15_25 = _RAND_1961[7:0];
  _RAND_1962 = {1{`RANDOM}};
  frameBuffer_15_26 = _RAND_1962[7:0];
  _RAND_1963 = {1{`RANDOM}};
  frameBuffer_15_27 = _RAND_1963[7:0];
  _RAND_1964 = {1{`RANDOM}};
  frameBuffer_15_28 = _RAND_1964[7:0];
  _RAND_1965 = {1{`RANDOM}};
  frameBuffer_15_29 = _RAND_1965[7:0];
  _RAND_1966 = {1{`RANDOM}};
  frameBuffer_15_30 = _RAND_1966[7:0];
  _RAND_1967 = {1{`RANDOM}};
  frameBuffer_15_31 = _RAND_1967[7:0];
  _RAND_1968 = {1{`RANDOM}};
  frameBuffer_15_32 = _RAND_1968[7:0];
  _RAND_1969 = {1{`RANDOM}};
  frameBuffer_15_33 = _RAND_1969[7:0];
  _RAND_1970 = {1{`RANDOM}};
  frameBuffer_15_34 = _RAND_1970[7:0];
  _RAND_1971 = {1{`RANDOM}};
  frameBuffer_15_35 = _RAND_1971[7:0];
  _RAND_1972 = {1{`RANDOM}};
  frameBuffer_15_36 = _RAND_1972[7:0];
  _RAND_1973 = {1{`RANDOM}};
  frameBuffer_15_37 = _RAND_1973[7:0];
  _RAND_1974 = {1{`RANDOM}};
  frameBuffer_15_38 = _RAND_1974[7:0];
  _RAND_1975 = {1{`RANDOM}};
  frameBuffer_15_39 = _RAND_1975[7:0];
  _RAND_1976 = {1{`RANDOM}};
  frameBuffer_15_40 = _RAND_1976[7:0];
  _RAND_1977 = {1{`RANDOM}};
  frameBuffer_15_41 = _RAND_1977[7:0];
  _RAND_1978 = {1{`RANDOM}};
  frameBuffer_15_42 = _RAND_1978[7:0];
  _RAND_1979 = {1{`RANDOM}};
  frameBuffer_15_43 = _RAND_1979[7:0];
  _RAND_1980 = {1{`RANDOM}};
  frameBuffer_15_44 = _RAND_1980[7:0];
  _RAND_1981 = {1{`RANDOM}};
  frameBuffer_15_45 = _RAND_1981[7:0];
  _RAND_1982 = {1{`RANDOM}};
  frameBuffer_15_46 = _RAND_1982[7:0];
  _RAND_1983 = {1{`RANDOM}};
  frameBuffer_15_47 = _RAND_1983[7:0];
  _RAND_1984 = {1{`RANDOM}};
  frameBuffer_15_48 = _RAND_1984[7:0];
  _RAND_1985 = {1{`RANDOM}};
  frameBuffer_15_49 = _RAND_1985[7:0];
  _RAND_1986 = {1{`RANDOM}};
  frameBuffer_15_50 = _RAND_1986[7:0];
  _RAND_1987 = {1{`RANDOM}};
  frameBuffer_15_51 = _RAND_1987[7:0];
  _RAND_1988 = {1{`RANDOM}};
  frameBuffer_15_52 = _RAND_1988[7:0];
  _RAND_1989 = {1{`RANDOM}};
  frameBuffer_15_53 = _RAND_1989[7:0];
  _RAND_1990 = {1{`RANDOM}};
  frameBuffer_15_54 = _RAND_1990[7:0];
  _RAND_1991 = {1{`RANDOM}};
  frameBuffer_15_55 = _RAND_1991[7:0];
  _RAND_1992 = {1{`RANDOM}};
  frameBuffer_15_56 = _RAND_1992[7:0];
  _RAND_1993 = {1{`RANDOM}};
  frameBuffer_15_57 = _RAND_1993[7:0];
  _RAND_1994 = {1{`RANDOM}};
  frameBuffer_15_58 = _RAND_1994[7:0];
  _RAND_1995 = {1{`RANDOM}};
  frameBuffer_15_59 = _RAND_1995[7:0];
  _RAND_1996 = {1{`RANDOM}};
  frameBuffer_15_60 = _RAND_1996[7:0];
  _RAND_1997 = {1{`RANDOM}};
  frameBuffer_15_61 = _RAND_1997[7:0];
  _RAND_1998 = {1{`RANDOM}};
  frameBuffer_15_62 = _RAND_1998[7:0];
  _RAND_1999 = {1{`RANDOM}};
  frameBuffer_15_63 = _RAND_1999[7:0];
  _RAND_2000 = {1{`RANDOM}};
  frameBuffer_15_64 = _RAND_2000[7:0];
  _RAND_2001 = {1{`RANDOM}};
  frameBuffer_15_65 = _RAND_2001[7:0];
  _RAND_2002 = {1{`RANDOM}};
  frameBuffer_15_66 = _RAND_2002[7:0];
  _RAND_2003 = {1{`RANDOM}};
  frameBuffer_15_67 = _RAND_2003[7:0];
  _RAND_2004 = {1{`RANDOM}};
  frameBuffer_15_68 = _RAND_2004[7:0];
  _RAND_2005 = {1{`RANDOM}};
  frameBuffer_15_69 = _RAND_2005[7:0];
  _RAND_2006 = {1{`RANDOM}};
  frameBuffer_15_70 = _RAND_2006[7:0];
  _RAND_2007 = {1{`RANDOM}};
  frameBuffer_15_71 = _RAND_2007[7:0];
  _RAND_2008 = {1{`RANDOM}};
  frameBuffer_15_72 = _RAND_2008[7:0];
  _RAND_2009 = {1{`RANDOM}};
  frameBuffer_15_73 = _RAND_2009[7:0];
  _RAND_2010 = {1{`RANDOM}};
  frameBuffer_15_74 = _RAND_2010[7:0];
  _RAND_2011 = {1{`RANDOM}};
  frameBuffer_15_75 = _RAND_2011[7:0];
  _RAND_2012 = {1{`RANDOM}};
  frameBuffer_15_76 = _RAND_2012[7:0];
  _RAND_2013 = {1{`RANDOM}};
  frameBuffer_15_77 = _RAND_2013[7:0];
  _RAND_2014 = {1{`RANDOM}};
  frameBuffer_15_78 = _RAND_2014[7:0];
  _RAND_2015 = {1{`RANDOM}};
  frameBuffer_15_79 = _RAND_2015[7:0];
  _RAND_2016 = {1{`RANDOM}};
  frameBuffer_15_80 = _RAND_2016[7:0];
  _RAND_2017 = {1{`RANDOM}};
  frameBuffer_15_81 = _RAND_2017[7:0];
  _RAND_2018 = {1{`RANDOM}};
  frameBuffer_15_82 = _RAND_2018[7:0];
  _RAND_2019 = {1{`RANDOM}};
  frameBuffer_15_83 = _RAND_2019[7:0];
  _RAND_2020 = {1{`RANDOM}};
  frameBuffer_15_84 = _RAND_2020[7:0];
  _RAND_2021 = {1{`RANDOM}};
  frameBuffer_15_85 = _RAND_2021[7:0];
  _RAND_2022 = {1{`RANDOM}};
  frameBuffer_15_86 = _RAND_2022[7:0];
  _RAND_2023 = {1{`RANDOM}};
  frameBuffer_15_87 = _RAND_2023[7:0];
  _RAND_2024 = {1{`RANDOM}};
  frameBuffer_15_88 = _RAND_2024[7:0];
  _RAND_2025 = {1{`RANDOM}};
  frameBuffer_15_89 = _RAND_2025[7:0];
  _RAND_2026 = {1{`RANDOM}};
  frameBuffer_15_90 = _RAND_2026[7:0];
  _RAND_2027 = {1{`RANDOM}};
  frameBuffer_15_91 = _RAND_2027[7:0];
  _RAND_2028 = {1{`RANDOM}};
  frameBuffer_15_92 = _RAND_2028[7:0];
  _RAND_2029 = {1{`RANDOM}};
  frameBuffer_15_93 = _RAND_2029[7:0];
  _RAND_2030 = {1{`RANDOM}};
  frameBuffer_15_94 = _RAND_2030[7:0];
  _RAND_2031 = {1{`RANDOM}};
  frameBuffer_15_95 = _RAND_2031[7:0];
  _RAND_2032 = {1{`RANDOM}};
  frameBuffer_15_96 = _RAND_2032[7:0];
  _RAND_2033 = {1{`RANDOM}};
  frameBuffer_15_97 = _RAND_2033[7:0];
  _RAND_2034 = {1{`RANDOM}};
  frameBuffer_15_98 = _RAND_2034[7:0];
  _RAND_2035 = {1{`RANDOM}};
  frameBuffer_15_99 = _RAND_2035[7:0];
  _RAND_2036 = {1{`RANDOM}};
  frameBuffer_15_100 = _RAND_2036[7:0];
  _RAND_2037 = {1{`RANDOM}};
  frameBuffer_15_101 = _RAND_2037[7:0];
  _RAND_2038 = {1{`RANDOM}};
  frameBuffer_15_102 = _RAND_2038[7:0];
  _RAND_2039 = {1{`RANDOM}};
  frameBuffer_15_103 = _RAND_2039[7:0];
  _RAND_2040 = {1{`RANDOM}};
  frameBuffer_15_104 = _RAND_2040[7:0];
  _RAND_2041 = {1{`RANDOM}};
  frameBuffer_15_105 = _RAND_2041[7:0];
  _RAND_2042 = {1{`RANDOM}};
  frameBuffer_15_106 = _RAND_2042[7:0];
  _RAND_2043 = {1{`RANDOM}};
  frameBuffer_15_107 = _RAND_2043[7:0];
  _RAND_2044 = {1{`RANDOM}};
  frameBuffer_15_108 = _RAND_2044[7:0];
  _RAND_2045 = {1{`RANDOM}};
  frameBuffer_15_109 = _RAND_2045[7:0];
  _RAND_2046 = {1{`RANDOM}};
  frameBuffer_15_110 = _RAND_2046[7:0];
  _RAND_2047 = {1{`RANDOM}};
  frameBuffer_15_111 = _RAND_2047[7:0];
  _RAND_2048 = {1{`RANDOM}};
  frameBuffer_15_112 = _RAND_2048[7:0];
  _RAND_2049 = {1{`RANDOM}};
  frameBuffer_15_113 = _RAND_2049[7:0];
  _RAND_2050 = {1{`RANDOM}};
  frameBuffer_15_114 = _RAND_2050[7:0];
  _RAND_2051 = {1{`RANDOM}};
  frameBuffer_15_115 = _RAND_2051[7:0];
  _RAND_2052 = {1{`RANDOM}};
  frameBuffer_15_116 = _RAND_2052[7:0];
  _RAND_2053 = {1{`RANDOM}};
  frameBuffer_15_117 = _RAND_2053[7:0];
  _RAND_2054 = {1{`RANDOM}};
  frameBuffer_15_118 = _RAND_2054[7:0];
  _RAND_2055 = {1{`RANDOM}};
  frameBuffer_15_119 = _RAND_2055[7:0];
  _RAND_2056 = {1{`RANDOM}};
  frameBuffer_15_120 = _RAND_2056[7:0];
  _RAND_2057 = {1{`RANDOM}};
  frameBuffer_15_121 = _RAND_2057[7:0];
  _RAND_2058 = {1{`RANDOM}};
  frameBuffer_15_122 = _RAND_2058[7:0];
  _RAND_2059 = {1{`RANDOM}};
  frameBuffer_15_123 = _RAND_2059[7:0];
  _RAND_2060 = {1{`RANDOM}};
  frameBuffer_15_124 = _RAND_2060[7:0];
  _RAND_2061 = {1{`RANDOM}};
  frameBuffer_15_125 = _RAND_2061[7:0];
  _RAND_2062 = {1{`RANDOM}};
  frameBuffer_15_126 = _RAND_2062[7:0];
  _RAND_2063 = {1{`RANDOM}};
  frameBuffer_15_127 = _RAND_2063[7:0];
  _RAND_2064 = {1{`RANDOM}};
  lineCounter = _RAND_2064[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
